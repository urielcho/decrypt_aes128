magic
tech sky130A
magscale 1 2
timestamp 1671591995
<< obsli1 >>
rect 1104 2159 358892 357425
<< obsm1 >>
rect 14 1912 359430 357456
<< metal2 >>
rect 18 359200 74 359800
rect 3882 359200 3938 359800
rect 7102 359200 7158 359800
rect 10966 359200 11022 359800
rect 14186 359200 14242 359800
rect 18050 359200 18106 359800
rect 21914 359200 21970 359800
rect 25134 359200 25190 359800
rect 28998 359200 29054 359800
rect 32862 359200 32918 359800
rect 36082 359200 36138 359800
rect 39946 359200 40002 359800
rect 43810 359200 43866 359800
rect 47030 359200 47086 359800
rect 50894 359200 50950 359800
rect 54758 359200 54814 359800
rect 57978 359200 58034 359800
rect 61842 359200 61898 359800
rect 65062 359200 65118 359800
rect 68926 359200 68982 359800
rect 72790 359200 72846 359800
rect 76010 359200 76066 359800
rect 79874 359200 79930 359800
rect 83738 359200 83794 359800
rect 86958 359200 87014 359800
rect 90822 359200 90878 359800
rect 94686 359200 94742 359800
rect 97906 359200 97962 359800
rect 101770 359200 101826 359800
rect 105634 359200 105690 359800
rect 108854 359200 108910 359800
rect 112718 359200 112774 359800
rect 115938 359200 115994 359800
rect 119802 359200 119858 359800
rect 123666 359200 123722 359800
rect 126886 359200 126942 359800
rect 130750 359200 130806 359800
rect 134614 359200 134670 359800
rect 137834 359200 137890 359800
rect 141698 359200 141754 359800
rect 145562 359200 145618 359800
rect 148782 359200 148838 359800
rect 152646 359200 152702 359800
rect 156510 359200 156566 359800
rect 159730 359200 159786 359800
rect 163594 359200 163650 359800
rect 166814 359200 166870 359800
rect 170678 359200 170734 359800
rect 174542 359200 174598 359800
rect 177762 359200 177818 359800
rect 181626 359200 181682 359800
rect 185490 359200 185546 359800
rect 188710 359200 188766 359800
rect 192574 359200 192630 359800
rect 196438 359200 196494 359800
rect 199658 359200 199714 359800
rect 203522 359200 203578 359800
rect 207386 359200 207442 359800
rect 210606 359200 210662 359800
rect 214470 359200 214526 359800
rect 217690 359200 217746 359800
rect 221554 359200 221610 359800
rect 225418 359200 225474 359800
rect 228638 359200 228694 359800
rect 232502 359200 232558 359800
rect 236366 359200 236422 359800
rect 239586 359200 239642 359800
rect 243450 359200 243506 359800
rect 247314 359200 247370 359800
rect 250534 359200 250590 359800
rect 254398 359200 254454 359800
rect 258262 359200 258318 359800
rect 261482 359200 261538 359800
rect 265346 359200 265402 359800
rect 268566 359200 268622 359800
rect 272430 359200 272486 359800
rect 276294 359200 276350 359800
rect 279514 359200 279570 359800
rect 283378 359200 283434 359800
rect 287242 359200 287298 359800
rect 290462 359200 290518 359800
rect 294326 359200 294382 359800
rect 298190 359200 298246 359800
rect 301410 359200 301466 359800
rect 305274 359200 305330 359800
rect 309138 359200 309194 359800
rect 312358 359200 312414 359800
rect 316222 359200 316278 359800
rect 319442 359200 319498 359800
rect 323306 359200 323362 359800
rect 327170 359200 327226 359800
rect 330390 359200 330446 359800
rect 334254 359200 334310 359800
rect 338118 359200 338174 359800
rect 341338 359200 341394 359800
rect 345202 359200 345258 359800
rect 349066 359200 349122 359800
rect 352286 359200 352342 359800
rect 356150 359200 356206 359800
rect 359370 359200 359426 359800
rect 18 200 74 800
rect 3238 200 3294 800
rect 7102 200 7158 800
rect 10322 200 10378 800
rect 14186 200 14242 800
rect 18050 200 18106 800
rect 21270 200 21326 800
rect 25134 200 25190 800
rect 28998 200 29054 800
rect 32218 200 32274 800
rect 36082 200 36138 800
rect 39946 200 40002 800
rect 43166 200 43222 800
rect 47030 200 47086 800
rect 50250 200 50306 800
rect 54114 200 54170 800
rect 57978 200 58034 800
rect 61198 200 61254 800
rect 65062 200 65118 800
rect 68926 200 68982 800
rect 72146 200 72202 800
rect 76010 200 76066 800
rect 79874 200 79930 800
rect 83094 200 83150 800
rect 86958 200 87014 800
rect 90822 200 90878 800
rect 94042 200 94098 800
rect 97906 200 97962 800
rect 101126 200 101182 800
rect 104990 200 105046 800
rect 108854 200 108910 800
rect 112074 200 112130 800
rect 115938 200 115994 800
rect 119802 200 119858 800
rect 123022 200 123078 800
rect 126886 200 126942 800
rect 130750 200 130806 800
rect 133970 200 134026 800
rect 137834 200 137890 800
rect 141698 200 141754 800
rect 144918 200 144974 800
rect 148782 200 148838 800
rect 152002 200 152058 800
rect 155866 200 155922 800
rect 159730 200 159786 800
rect 162950 200 163006 800
rect 166814 200 166870 800
rect 170678 200 170734 800
rect 173898 200 173954 800
rect 177762 200 177818 800
rect 181626 200 181682 800
rect 184846 200 184902 800
rect 188710 200 188766 800
rect 192574 200 192630 800
rect 195794 200 195850 800
rect 199658 200 199714 800
rect 202878 200 202934 800
rect 206742 200 206798 800
rect 210606 200 210662 800
rect 213826 200 213882 800
rect 217690 200 217746 800
rect 221554 200 221610 800
rect 224774 200 224830 800
rect 228638 200 228694 800
rect 232502 200 232558 800
rect 235722 200 235778 800
rect 239586 200 239642 800
rect 243450 200 243506 800
rect 246670 200 246726 800
rect 250534 200 250590 800
rect 253754 200 253810 800
rect 257618 200 257674 800
rect 261482 200 261538 800
rect 264702 200 264758 800
rect 268566 200 268622 800
rect 272430 200 272486 800
rect 275650 200 275706 800
rect 279514 200 279570 800
rect 283378 200 283434 800
rect 286598 200 286654 800
rect 290462 200 290518 800
rect 294326 200 294382 800
rect 297546 200 297602 800
rect 301410 200 301466 800
rect 304630 200 304686 800
rect 308494 200 308550 800
rect 312358 200 312414 800
rect 315578 200 315634 800
rect 319442 200 319498 800
rect 323306 200 323362 800
rect 326526 200 326582 800
rect 330390 200 330446 800
rect 334254 200 334310 800
rect 337474 200 337530 800
rect 341338 200 341394 800
rect 345202 200 345258 800
rect 348422 200 348478 800
rect 352286 200 352342 800
rect 355506 200 355562 800
rect 359370 200 359426 800
<< obsm2 >>
rect 130 359144 3826 359258
rect 3994 359144 7046 359258
rect 7214 359144 10910 359258
rect 11078 359144 14130 359258
rect 14298 359144 17994 359258
rect 18162 359144 21858 359258
rect 22026 359144 25078 359258
rect 25246 359144 28942 359258
rect 29110 359144 32806 359258
rect 32974 359144 36026 359258
rect 36194 359144 39890 359258
rect 40058 359144 43754 359258
rect 43922 359144 46974 359258
rect 47142 359144 50838 359258
rect 51006 359144 54702 359258
rect 54870 359144 57922 359258
rect 58090 359144 61786 359258
rect 61954 359144 65006 359258
rect 65174 359144 68870 359258
rect 69038 359144 72734 359258
rect 72902 359144 75954 359258
rect 76122 359144 79818 359258
rect 79986 359144 83682 359258
rect 83850 359144 86902 359258
rect 87070 359144 90766 359258
rect 90934 359144 94630 359258
rect 94798 359144 97850 359258
rect 98018 359144 101714 359258
rect 101882 359144 105578 359258
rect 105746 359144 108798 359258
rect 108966 359144 112662 359258
rect 112830 359144 115882 359258
rect 116050 359144 119746 359258
rect 119914 359144 123610 359258
rect 123778 359144 126830 359258
rect 126998 359144 130694 359258
rect 130862 359144 134558 359258
rect 134726 359144 137778 359258
rect 137946 359144 141642 359258
rect 141810 359144 145506 359258
rect 145674 359144 148726 359258
rect 148894 359144 152590 359258
rect 152758 359144 156454 359258
rect 156622 359144 159674 359258
rect 159842 359144 163538 359258
rect 163706 359144 166758 359258
rect 166926 359144 170622 359258
rect 170790 359144 174486 359258
rect 174654 359144 177706 359258
rect 177874 359144 181570 359258
rect 181738 359144 185434 359258
rect 185602 359144 188654 359258
rect 188822 359144 192518 359258
rect 192686 359144 196382 359258
rect 196550 359144 199602 359258
rect 199770 359144 203466 359258
rect 203634 359144 207330 359258
rect 207498 359144 210550 359258
rect 210718 359144 214414 359258
rect 214582 359144 217634 359258
rect 217802 359144 221498 359258
rect 221666 359144 225362 359258
rect 225530 359144 228582 359258
rect 228750 359144 232446 359258
rect 232614 359144 236310 359258
rect 236478 359144 239530 359258
rect 239698 359144 243394 359258
rect 243562 359144 247258 359258
rect 247426 359144 250478 359258
rect 250646 359144 254342 359258
rect 254510 359144 258206 359258
rect 258374 359144 261426 359258
rect 261594 359144 265290 359258
rect 265458 359144 268510 359258
rect 268678 359144 272374 359258
rect 272542 359144 276238 359258
rect 276406 359144 279458 359258
rect 279626 359144 283322 359258
rect 283490 359144 287186 359258
rect 287354 359144 290406 359258
rect 290574 359144 294270 359258
rect 294438 359144 298134 359258
rect 298302 359144 301354 359258
rect 301522 359144 305218 359258
rect 305386 359144 309082 359258
rect 309250 359144 312302 359258
rect 312470 359144 316166 359258
rect 316334 359144 319386 359258
rect 319554 359144 323250 359258
rect 323418 359144 327114 359258
rect 327282 359144 330334 359258
rect 330502 359144 334198 359258
rect 334366 359144 338062 359258
rect 338230 359144 341282 359258
rect 341450 359144 345146 359258
rect 345314 359144 349010 359258
rect 349178 359144 352230 359258
rect 352398 359144 356094 359258
rect 356262 359144 359314 359258
rect 20 856 359424 359144
rect 130 734 3182 856
rect 3350 734 7046 856
rect 7214 734 10266 856
rect 10434 734 14130 856
rect 14298 734 17994 856
rect 18162 734 21214 856
rect 21382 734 25078 856
rect 25246 734 28942 856
rect 29110 734 32162 856
rect 32330 734 36026 856
rect 36194 734 39890 856
rect 40058 734 43110 856
rect 43278 734 46974 856
rect 47142 734 50194 856
rect 50362 734 54058 856
rect 54226 734 57922 856
rect 58090 734 61142 856
rect 61310 734 65006 856
rect 65174 734 68870 856
rect 69038 734 72090 856
rect 72258 734 75954 856
rect 76122 734 79818 856
rect 79986 734 83038 856
rect 83206 734 86902 856
rect 87070 734 90766 856
rect 90934 734 93986 856
rect 94154 734 97850 856
rect 98018 734 101070 856
rect 101238 734 104934 856
rect 105102 734 108798 856
rect 108966 734 112018 856
rect 112186 734 115882 856
rect 116050 734 119746 856
rect 119914 734 122966 856
rect 123134 734 126830 856
rect 126998 734 130694 856
rect 130862 734 133914 856
rect 134082 734 137778 856
rect 137946 734 141642 856
rect 141810 734 144862 856
rect 145030 734 148726 856
rect 148894 734 151946 856
rect 152114 734 155810 856
rect 155978 734 159674 856
rect 159842 734 162894 856
rect 163062 734 166758 856
rect 166926 734 170622 856
rect 170790 734 173842 856
rect 174010 734 177706 856
rect 177874 734 181570 856
rect 181738 734 184790 856
rect 184958 734 188654 856
rect 188822 734 192518 856
rect 192686 734 195738 856
rect 195906 734 199602 856
rect 199770 734 202822 856
rect 202990 734 206686 856
rect 206854 734 210550 856
rect 210718 734 213770 856
rect 213938 734 217634 856
rect 217802 734 221498 856
rect 221666 734 224718 856
rect 224886 734 228582 856
rect 228750 734 232446 856
rect 232614 734 235666 856
rect 235834 734 239530 856
rect 239698 734 243394 856
rect 243562 734 246614 856
rect 246782 734 250478 856
rect 250646 734 253698 856
rect 253866 734 257562 856
rect 257730 734 261426 856
rect 261594 734 264646 856
rect 264814 734 268510 856
rect 268678 734 272374 856
rect 272542 734 275594 856
rect 275762 734 279458 856
rect 279626 734 283322 856
rect 283490 734 286542 856
rect 286710 734 290406 856
rect 290574 734 294270 856
rect 294438 734 297490 856
rect 297658 734 301354 856
rect 301522 734 304574 856
rect 304742 734 308438 856
rect 308606 734 312302 856
rect 312470 734 315522 856
rect 315690 734 319386 856
rect 319554 734 323250 856
rect 323418 734 326470 856
rect 326638 734 330334 856
rect 330502 734 334198 856
rect 334366 734 337418 856
rect 337586 734 341282 856
rect 341450 734 345146 856
rect 345314 734 348366 856
rect 348534 734 352230 856
rect 352398 734 355450 856
rect 355618 734 359314 856
<< metal3 >>
rect 200 356328 800 356448
rect 359200 356328 359800 356448
rect 200 352928 800 353048
rect 359200 352248 359800 352368
rect 200 348848 800 348968
rect 359200 348848 359800 348968
rect 200 344768 800 344888
rect 359200 344768 359800 344888
rect 200 341368 800 341488
rect 359200 340688 359800 340808
rect 200 337288 800 337408
rect 359200 337288 359800 337408
rect 200 333208 800 333328
rect 359200 333208 359800 333328
rect 200 329808 800 329928
rect 359200 329128 359800 329248
rect 200 325728 800 325848
rect 359200 325728 359800 325848
rect 200 321648 800 321768
rect 359200 321648 359800 321768
rect 200 318248 800 318368
rect 359200 317568 359800 317688
rect 200 314168 800 314288
rect 359200 314168 359800 314288
rect 200 310768 800 310888
rect 359200 310088 359800 310208
rect 200 306688 800 306808
rect 359200 306688 359800 306808
rect 200 302608 800 302728
rect 359200 302608 359800 302728
rect 200 299208 800 299328
rect 359200 298528 359800 298648
rect 200 295128 800 295248
rect 359200 295128 359800 295248
rect 200 291048 800 291168
rect 359200 291048 359800 291168
rect 200 287648 800 287768
rect 359200 286968 359800 287088
rect 200 283568 800 283688
rect 359200 283568 359800 283688
rect 200 279488 800 279608
rect 359200 279488 359800 279608
rect 200 276088 800 276208
rect 359200 275408 359800 275528
rect 200 272008 800 272128
rect 359200 272008 359800 272128
rect 200 267928 800 268048
rect 359200 267928 359800 268048
rect 200 264528 800 264648
rect 359200 263848 359800 263968
rect 200 260448 800 260568
rect 359200 260448 359800 260568
rect 200 257048 800 257168
rect 359200 256368 359800 256488
rect 200 252968 800 253088
rect 359200 252968 359800 253088
rect 200 248888 800 249008
rect 359200 248888 359800 249008
rect 200 245488 800 245608
rect 359200 244808 359800 244928
rect 200 241408 800 241528
rect 359200 241408 359800 241528
rect 200 237328 800 237448
rect 359200 237328 359800 237448
rect 200 233928 800 234048
rect 359200 233248 359800 233368
rect 200 229848 800 229968
rect 359200 229848 359800 229968
rect 200 225768 800 225888
rect 359200 225768 359800 225888
rect 200 222368 800 222488
rect 359200 221688 359800 221808
rect 200 218288 800 218408
rect 359200 218288 359800 218408
rect 200 214208 800 214328
rect 359200 214208 359800 214328
rect 200 210808 800 210928
rect 359200 210128 359800 210248
rect 200 206728 800 206848
rect 359200 206728 359800 206848
rect 200 203328 800 203448
rect 359200 202648 359800 202768
rect 200 199248 800 199368
rect 359200 199248 359800 199368
rect 200 195168 800 195288
rect 359200 195168 359800 195288
rect 200 191768 800 191888
rect 359200 191088 359800 191208
rect 200 187688 800 187808
rect 359200 187688 359800 187808
rect 200 183608 800 183728
rect 359200 183608 359800 183728
rect 200 180208 800 180328
rect 359200 179528 359800 179648
rect 200 176128 800 176248
rect 359200 176128 359800 176248
rect 200 172048 800 172168
rect 359200 172048 359800 172168
rect 200 168648 800 168768
rect 359200 167968 359800 168088
rect 200 164568 800 164688
rect 359200 164568 359800 164688
rect 200 160488 800 160608
rect 359200 160488 359800 160608
rect 200 157088 800 157208
rect 359200 156408 359800 156528
rect 200 153008 800 153128
rect 359200 153008 359800 153128
rect 200 149608 800 149728
rect 359200 148928 359800 149048
rect 200 145528 800 145648
rect 359200 145528 359800 145648
rect 200 141448 800 141568
rect 359200 141448 359800 141568
rect 200 138048 800 138168
rect 359200 137368 359800 137488
rect 200 133968 800 134088
rect 359200 133968 359800 134088
rect 200 129888 800 130008
rect 359200 129888 359800 130008
rect 200 126488 800 126608
rect 359200 125808 359800 125928
rect 200 122408 800 122528
rect 359200 122408 359800 122528
rect 200 118328 800 118448
rect 359200 118328 359800 118448
rect 200 114928 800 115048
rect 359200 114248 359800 114368
rect 200 110848 800 110968
rect 359200 110848 359800 110968
rect 200 106768 800 106888
rect 359200 106768 359800 106888
rect 200 103368 800 103488
rect 359200 102688 359800 102808
rect 200 99288 800 99408
rect 359200 99288 359800 99408
rect 200 95888 800 96008
rect 359200 95208 359800 95328
rect 200 91808 800 91928
rect 359200 91808 359800 91928
rect 200 87728 800 87848
rect 359200 87728 359800 87848
rect 200 84328 800 84448
rect 359200 83648 359800 83768
rect 200 80248 800 80368
rect 359200 80248 359800 80368
rect 200 76168 800 76288
rect 359200 76168 359800 76288
rect 200 72768 800 72888
rect 359200 72088 359800 72208
rect 200 68688 800 68808
rect 359200 68688 359800 68808
rect 200 64608 800 64728
rect 359200 64608 359800 64728
rect 200 61208 800 61328
rect 359200 60528 359800 60648
rect 200 57128 800 57248
rect 359200 57128 359800 57248
rect 200 53048 800 53168
rect 359200 53048 359800 53168
rect 200 49648 800 49768
rect 359200 48968 359800 49088
rect 200 45568 800 45688
rect 359200 45568 359800 45688
rect 200 42168 800 42288
rect 359200 41488 359800 41608
rect 200 38088 800 38208
rect 359200 38088 359800 38208
rect 200 34008 800 34128
rect 359200 34008 359800 34128
rect 200 30608 800 30728
rect 359200 29928 359800 30048
rect 200 26528 800 26648
rect 359200 26528 359800 26648
rect 200 22448 800 22568
rect 359200 22448 359800 22568
rect 200 19048 800 19168
rect 359200 18368 359800 18488
rect 200 14968 800 15088
rect 359200 14968 359800 15088
rect 200 10888 800 11008
rect 359200 10888 359800 11008
rect 200 7488 800 7608
rect 359200 6808 359800 6928
rect 200 3408 800 3528
rect 359200 3408 359800 3528
<< obsm3 >>
rect 800 356528 359200 357441
rect 880 356248 359120 356528
rect 800 353128 359200 356248
rect 880 352848 359200 353128
rect 800 352448 359200 352848
rect 800 352168 359120 352448
rect 800 349048 359200 352168
rect 880 348768 359120 349048
rect 800 344968 359200 348768
rect 880 344688 359120 344968
rect 800 341568 359200 344688
rect 880 341288 359200 341568
rect 800 340888 359200 341288
rect 800 340608 359120 340888
rect 800 337488 359200 340608
rect 880 337208 359120 337488
rect 800 333408 359200 337208
rect 880 333128 359120 333408
rect 800 330008 359200 333128
rect 880 329728 359200 330008
rect 800 329328 359200 329728
rect 800 329048 359120 329328
rect 800 325928 359200 329048
rect 880 325648 359120 325928
rect 800 321848 359200 325648
rect 880 321568 359120 321848
rect 800 318448 359200 321568
rect 880 318168 359200 318448
rect 800 317768 359200 318168
rect 800 317488 359120 317768
rect 800 314368 359200 317488
rect 880 314088 359120 314368
rect 800 310968 359200 314088
rect 880 310688 359200 310968
rect 800 310288 359200 310688
rect 800 310008 359120 310288
rect 800 306888 359200 310008
rect 880 306608 359120 306888
rect 800 302808 359200 306608
rect 880 302528 359120 302808
rect 800 299408 359200 302528
rect 880 299128 359200 299408
rect 800 298728 359200 299128
rect 800 298448 359120 298728
rect 800 295328 359200 298448
rect 880 295048 359120 295328
rect 800 291248 359200 295048
rect 880 290968 359120 291248
rect 800 287848 359200 290968
rect 880 287568 359200 287848
rect 800 287168 359200 287568
rect 800 286888 359120 287168
rect 800 283768 359200 286888
rect 880 283488 359120 283768
rect 800 279688 359200 283488
rect 880 279408 359120 279688
rect 800 276288 359200 279408
rect 880 276008 359200 276288
rect 800 275608 359200 276008
rect 800 275328 359120 275608
rect 800 272208 359200 275328
rect 880 271928 359120 272208
rect 800 268128 359200 271928
rect 880 267848 359120 268128
rect 800 264728 359200 267848
rect 880 264448 359200 264728
rect 800 264048 359200 264448
rect 800 263768 359120 264048
rect 800 260648 359200 263768
rect 880 260368 359120 260648
rect 800 257248 359200 260368
rect 880 256968 359200 257248
rect 800 256568 359200 256968
rect 800 256288 359120 256568
rect 800 253168 359200 256288
rect 880 252888 359120 253168
rect 800 249088 359200 252888
rect 880 248808 359120 249088
rect 800 245688 359200 248808
rect 880 245408 359200 245688
rect 800 245008 359200 245408
rect 800 244728 359120 245008
rect 800 241608 359200 244728
rect 880 241328 359120 241608
rect 800 237528 359200 241328
rect 880 237248 359120 237528
rect 800 234128 359200 237248
rect 880 233848 359200 234128
rect 800 233448 359200 233848
rect 800 233168 359120 233448
rect 800 230048 359200 233168
rect 880 229768 359120 230048
rect 800 225968 359200 229768
rect 880 225688 359120 225968
rect 800 222568 359200 225688
rect 880 222288 359200 222568
rect 800 221888 359200 222288
rect 800 221608 359120 221888
rect 800 218488 359200 221608
rect 880 218208 359120 218488
rect 800 214408 359200 218208
rect 880 214128 359120 214408
rect 800 211008 359200 214128
rect 880 210728 359200 211008
rect 800 210328 359200 210728
rect 800 210048 359120 210328
rect 800 206928 359200 210048
rect 880 206648 359120 206928
rect 800 203528 359200 206648
rect 880 203248 359200 203528
rect 800 202848 359200 203248
rect 800 202568 359120 202848
rect 800 199448 359200 202568
rect 880 199168 359120 199448
rect 800 195368 359200 199168
rect 880 195088 359120 195368
rect 800 191968 359200 195088
rect 880 191688 359200 191968
rect 800 191288 359200 191688
rect 800 191008 359120 191288
rect 800 187888 359200 191008
rect 880 187608 359120 187888
rect 800 183808 359200 187608
rect 880 183528 359120 183808
rect 800 180408 359200 183528
rect 880 180128 359200 180408
rect 800 179728 359200 180128
rect 800 179448 359120 179728
rect 800 176328 359200 179448
rect 880 176048 359120 176328
rect 800 172248 359200 176048
rect 880 171968 359120 172248
rect 800 168848 359200 171968
rect 880 168568 359200 168848
rect 800 168168 359200 168568
rect 800 167888 359120 168168
rect 800 164768 359200 167888
rect 880 164488 359120 164768
rect 800 160688 359200 164488
rect 880 160408 359120 160688
rect 800 157288 359200 160408
rect 880 157008 359200 157288
rect 800 156608 359200 157008
rect 800 156328 359120 156608
rect 800 153208 359200 156328
rect 880 152928 359120 153208
rect 800 149808 359200 152928
rect 880 149528 359200 149808
rect 800 149128 359200 149528
rect 800 148848 359120 149128
rect 800 145728 359200 148848
rect 880 145448 359120 145728
rect 800 141648 359200 145448
rect 880 141368 359120 141648
rect 800 138248 359200 141368
rect 880 137968 359200 138248
rect 800 137568 359200 137968
rect 800 137288 359120 137568
rect 800 134168 359200 137288
rect 880 133888 359120 134168
rect 800 130088 359200 133888
rect 880 129808 359120 130088
rect 800 126688 359200 129808
rect 880 126408 359200 126688
rect 800 126008 359200 126408
rect 800 125728 359120 126008
rect 800 122608 359200 125728
rect 880 122328 359120 122608
rect 800 118528 359200 122328
rect 880 118248 359120 118528
rect 800 115128 359200 118248
rect 880 114848 359200 115128
rect 800 114448 359200 114848
rect 800 114168 359120 114448
rect 800 111048 359200 114168
rect 880 110768 359120 111048
rect 800 106968 359200 110768
rect 880 106688 359120 106968
rect 800 103568 359200 106688
rect 880 103288 359200 103568
rect 800 102888 359200 103288
rect 800 102608 359120 102888
rect 800 99488 359200 102608
rect 880 99208 359120 99488
rect 800 96088 359200 99208
rect 880 95808 359200 96088
rect 800 95408 359200 95808
rect 800 95128 359120 95408
rect 800 92008 359200 95128
rect 880 91728 359120 92008
rect 800 87928 359200 91728
rect 880 87648 359120 87928
rect 800 84528 359200 87648
rect 880 84248 359200 84528
rect 800 83848 359200 84248
rect 800 83568 359120 83848
rect 800 80448 359200 83568
rect 880 80168 359120 80448
rect 800 76368 359200 80168
rect 880 76088 359120 76368
rect 800 72968 359200 76088
rect 880 72688 359200 72968
rect 800 72288 359200 72688
rect 800 72008 359120 72288
rect 800 68888 359200 72008
rect 880 68608 359120 68888
rect 800 64808 359200 68608
rect 880 64528 359120 64808
rect 800 61408 359200 64528
rect 880 61128 359200 61408
rect 800 60728 359200 61128
rect 800 60448 359120 60728
rect 800 57328 359200 60448
rect 880 57048 359120 57328
rect 800 53248 359200 57048
rect 880 52968 359120 53248
rect 800 49848 359200 52968
rect 880 49568 359200 49848
rect 800 49168 359200 49568
rect 800 48888 359120 49168
rect 800 45768 359200 48888
rect 880 45488 359120 45768
rect 800 42368 359200 45488
rect 880 42088 359200 42368
rect 800 41688 359200 42088
rect 800 41408 359120 41688
rect 800 38288 359200 41408
rect 880 38008 359120 38288
rect 800 34208 359200 38008
rect 880 33928 359120 34208
rect 800 30808 359200 33928
rect 880 30528 359200 30808
rect 800 30128 359200 30528
rect 800 29848 359120 30128
rect 800 26728 359200 29848
rect 880 26448 359120 26728
rect 800 22648 359200 26448
rect 880 22368 359120 22648
rect 800 19248 359200 22368
rect 880 18968 359200 19248
rect 800 18568 359200 18968
rect 800 18288 359120 18568
rect 800 15168 359200 18288
rect 880 14888 359120 15168
rect 800 11088 359200 14888
rect 880 10808 359120 11088
rect 800 7688 359200 10808
rect 880 7408 359200 7688
rect 800 7008 359200 7408
rect 800 6728 359120 7008
rect 800 3608 359200 6728
rect 880 3328 359120 3608
rect 800 1531 359200 3328
<< metal4 >>
rect 4208 2128 4528 357456
rect 19568 2128 19888 357456
rect 34928 2128 35248 357456
rect 50288 2128 50608 357456
rect 65648 2128 65968 357456
rect 81008 2128 81328 357456
rect 96368 2128 96688 357456
rect 111728 2128 112048 357456
rect 127088 2128 127408 357456
rect 142448 2128 142768 357456
rect 157808 2128 158128 357456
rect 173168 2128 173488 357456
rect 188528 2128 188848 357456
rect 203888 2128 204208 357456
rect 219248 2128 219568 357456
rect 234608 2128 234928 357456
rect 249968 2128 250288 357456
rect 265328 2128 265648 357456
rect 280688 2128 281008 357456
rect 296048 2128 296368 357456
rect 311408 2128 311728 357456
rect 326768 2128 327088 357456
rect 342128 2128 342448 357456
rect 357488 2128 357808 357456
<< obsm4 >>
rect 6315 2048 19488 357237
rect 19968 2048 34848 357237
rect 35328 2048 50208 357237
rect 50688 2048 65568 357237
rect 66048 2048 80928 357237
rect 81408 2048 96288 357237
rect 96768 2048 111648 357237
rect 112128 2048 127008 357237
rect 127488 2048 142368 357237
rect 142848 2048 157728 357237
rect 158208 2048 173088 357237
rect 173568 2048 188448 357237
rect 188928 2048 203808 357237
rect 204288 2048 219168 357237
rect 219648 2048 234528 357237
rect 235008 2048 249888 357237
rect 250368 2048 265248 357237
rect 265728 2048 280608 357237
rect 281088 2048 295968 357237
rect 296448 2048 311328 357237
rect 311808 2048 326688 357237
rect 327168 2048 342048 357237
rect 342528 2048 353773 357237
rect 6315 1531 353773 2048
<< labels >>
rlabel metal3 s 359200 298528 359800 298648 6 clk
port 1 nsew signal input
rlabel metal2 s 341338 200 341394 800 6 decReset
port 2 nsew signal input
rlabel metal3 s 359200 34008 359800 34128 6 in[0]
port 3 nsew signal input
rlabel metal3 s 200 333208 800 333328 6 in[100]
port 4 nsew signal input
rlabel metal3 s 200 337288 800 337408 6 in[101]
port 5 nsew signal input
rlabel metal2 s 290462 200 290518 800 6 in[102]
port 6 nsew signal input
rlabel metal3 s 359200 72088 359800 72208 6 in[103]
port 7 nsew signal input
rlabel metal2 s 185490 359200 185546 359800 6 in[104]
port 8 nsew signal input
rlabel metal3 s 200 30608 800 30728 6 in[105]
port 9 nsew signal input
rlabel metal3 s 200 241408 800 241528 6 in[106]
port 10 nsew signal input
rlabel metal2 s 148782 359200 148838 359800 6 in[107]
port 11 nsew signal input
rlabel metal2 s 214470 359200 214526 359800 6 in[108]
port 12 nsew signal input
rlabel metal2 s 247314 359200 247370 359800 6 in[109]
port 13 nsew signal input
rlabel metal2 s 86958 359200 87014 359800 6 in[10]
port 14 nsew signal input
rlabel metal2 s 319442 359200 319498 359800 6 in[110]
port 15 nsew signal input
rlabel metal3 s 200 95888 800 96008 6 in[111]
port 16 nsew signal input
rlabel metal2 s 352286 200 352342 800 6 in[112]
port 17 nsew signal input
rlabel metal2 s 79874 200 79930 800 6 in[113]
port 18 nsew signal input
rlabel metal3 s 200 210808 800 210928 6 in[114]
port 19 nsew signal input
rlabel metal3 s 200 203328 800 203448 6 in[115]
port 20 nsew signal input
rlabel metal2 s 268566 359200 268622 359800 6 in[116]
port 21 nsew signal input
rlabel metal3 s 359200 340688 359800 340808 6 in[117]
port 22 nsew signal input
rlabel metal2 s 65062 359200 65118 359800 6 in[118]
port 23 nsew signal input
rlabel metal3 s 359200 102688 359800 102808 6 in[119]
port 24 nsew signal input
rlabel metal3 s 200 295128 800 295248 6 in[11]
port 25 nsew signal input
rlabel metal3 s 359200 221688 359800 221808 6 in[120]
port 26 nsew signal input
rlabel metal2 s 272430 200 272486 800 6 in[121]
port 27 nsew signal input
rlabel metal2 s 130750 200 130806 800 6 in[122]
port 28 nsew signal input
rlabel metal2 s 119802 359200 119858 359800 6 in[123]
port 29 nsew signal input
rlabel metal3 s 359200 179528 359800 179648 6 in[124]
port 30 nsew signal input
rlabel metal2 s 246670 200 246726 800 6 in[125]
port 31 nsew signal input
rlabel metal3 s 359200 260448 359800 260568 6 in[126]
port 32 nsew signal input
rlabel metal3 s 359200 267928 359800 268048 6 in[127]
port 33 nsew signal input
rlabel metal2 s 83094 200 83150 800 6 in[12]
port 34 nsew signal input
rlabel metal3 s 359200 187688 359800 187808 6 in[13]
port 35 nsew signal input
rlabel metal2 s 21270 200 21326 800 6 in[14]
port 36 nsew signal input
rlabel metal3 s 200 279488 800 279608 6 in[15]
port 37 nsew signal input
rlabel metal3 s 200 267928 800 268048 6 in[16]
port 38 nsew signal input
rlabel metal3 s 200 114928 800 115048 6 in[17]
port 39 nsew signal input
rlabel metal3 s 200 321648 800 321768 6 in[18]
port 40 nsew signal input
rlabel metal2 s 345202 359200 345258 359800 6 in[19]
port 41 nsew signal input
rlabel metal3 s 359200 110848 359800 110968 6 in[1]
port 42 nsew signal input
rlabel metal2 s 232502 200 232558 800 6 in[20]
port 43 nsew signal input
rlabel metal3 s 359200 241408 359800 241528 6 in[21]
port 44 nsew signal input
rlabel metal2 s 184846 200 184902 800 6 in[22]
port 45 nsew signal input
rlabel metal3 s 359200 356328 359800 356448 6 in[23]
port 46 nsew signal input
rlabel metal2 s 250534 359200 250590 359800 6 in[24]
port 47 nsew signal input
rlabel metal2 s 3882 359200 3938 359800 6 in[25]
port 48 nsew signal input
rlabel metal3 s 200 22448 800 22568 6 in[26]
port 49 nsew signal input
rlabel metal3 s 359200 141448 359800 141568 6 in[27]
port 50 nsew signal input
rlabel metal3 s 359200 87728 359800 87848 6 in[28]
port 51 nsew signal input
rlabel metal2 s 32218 200 32274 800 6 in[29]
port 52 nsew signal input
rlabel metal3 s 200 187688 800 187808 6 in[2]
port 53 nsew signal input
rlabel metal3 s 200 3408 800 3528 6 in[30]
port 54 nsew signal input
rlabel metal2 s 21914 359200 21970 359800 6 in[31]
port 55 nsew signal input
rlabel metal3 s 359200 306688 359800 306808 6 in[32]
port 56 nsew signal input
rlabel metal2 s 217690 359200 217746 359800 6 in[33]
port 57 nsew signal input
rlabel metal2 s 126886 359200 126942 359800 6 in[34]
port 58 nsew signal input
rlabel metal3 s 200 133968 800 134088 6 in[35]
port 59 nsew signal input
rlabel metal3 s 359200 80248 359800 80368 6 in[36]
port 60 nsew signal input
rlabel metal3 s 359200 156408 359800 156528 6 in[37]
port 61 nsew signal input
rlabel metal3 s 359200 183608 359800 183728 6 in[38]
port 62 nsew signal input
rlabel metal2 s 221554 200 221610 800 6 in[39]
port 63 nsew signal input
rlabel metal3 s 359200 76168 359800 76288 6 in[3]
port 64 nsew signal input
rlabel metal3 s 200 153008 800 153128 6 in[40]
port 65 nsew signal input
rlabel metal2 s 90822 359200 90878 359800 6 in[41]
port 66 nsew signal input
rlabel metal2 s 304630 200 304686 800 6 in[42]
port 67 nsew signal input
rlabel metal3 s 200 237328 800 237448 6 in[43]
port 68 nsew signal input
rlabel metal2 s 250534 200 250590 800 6 in[44]
port 69 nsew signal input
rlabel metal2 s 225418 359200 225474 359800 6 in[45]
port 70 nsew signal input
rlabel metal2 s 97906 359200 97962 359800 6 in[46]
port 71 nsew signal input
rlabel metal3 s 200 344768 800 344888 6 in[47]
port 72 nsew signal input
rlabel metal2 s 210606 359200 210662 359800 6 in[48]
port 73 nsew signal input
rlabel metal2 s 177762 200 177818 800 6 in[49]
port 74 nsew signal input
rlabel metal3 s 359200 41488 359800 41608 6 in[4]
port 75 nsew signal input
rlabel metal2 s 156510 359200 156566 359800 6 in[50]
port 76 nsew signal input
rlabel metal2 s 152002 200 152058 800 6 in[51]
port 77 nsew signal input
rlabel metal3 s 200 103368 800 103488 6 in[52]
port 78 nsew signal input
rlabel metal2 s 141698 359200 141754 359800 6 in[53]
port 79 nsew signal input
rlabel metal2 s 232502 359200 232558 359800 6 in[54]
port 80 nsew signal input
rlabel metal3 s 359200 291048 359800 291168 6 in[55]
port 81 nsew signal input
rlabel metal2 s 39946 200 40002 800 6 in[56]
port 82 nsew signal input
rlabel metal2 s 202878 200 202934 800 6 in[57]
port 83 nsew signal input
rlabel metal3 s 359200 337288 359800 337408 6 in[58]
port 84 nsew signal input
rlabel metal2 s 76010 359200 76066 359800 6 in[59]
port 85 nsew signal input
rlabel metal2 s 334254 359200 334310 359800 6 in[5]
port 86 nsew signal input
rlabel metal3 s 200 172048 800 172168 6 in[60]
port 87 nsew signal input
rlabel metal3 s 359200 295128 359800 295248 6 in[61]
port 88 nsew signal input
rlabel metal3 s 200 138048 800 138168 6 in[62]
port 89 nsew signal input
rlabel metal2 s 170678 359200 170734 359800 6 in[63]
port 90 nsew signal input
rlabel metal3 s 359200 60528 359800 60648 6 in[64]
port 91 nsew signal input
rlabel metal3 s 359200 125808 359800 125928 6 in[65]
port 92 nsew signal input
rlabel metal2 s 326526 200 326582 800 6 in[66]
port 93 nsew signal input
rlabel metal3 s 359200 314168 359800 314288 6 in[67]
port 94 nsew signal input
rlabel metal3 s 200 87728 800 87848 6 in[68]
port 95 nsew signal input
rlabel metal2 s 28998 359200 29054 359800 6 in[69]
port 96 nsew signal input
rlabel metal2 s 94686 359200 94742 359800 6 in[6]
port 97 nsew signal input
rlabel metal3 s 359200 26528 359800 26648 6 in[70]
port 98 nsew signal input
rlabel metal3 s 200 276088 800 276208 6 in[71]
port 99 nsew signal input
rlabel metal3 s 200 287648 800 287768 6 in[72]
port 100 nsew signal input
rlabel metal3 s 359200 286968 359800 287088 6 in[73]
port 101 nsew signal input
rlabel metal3 s 359200 164568 359800 164688 6 in[74]
port 102 nsew signal input
rlabel metal3 s 359200 283568 359800 283688 6 in[75]
port 103 nsew signal input
rlabel metal3 s 359200 244808 359800 244928 6 in[76]
port 104 nsew signal input
rlabel metal2 s 14186 359200 14242 359800 6 in[77]
port 105 nsew signal input
rlabel metal3 s 359200 10888 359800 11008 6 in[78]
port 106 nsew signal input
rlabel metal2 s 57978 359200 58034 359800 6 in[79]
port 107 nsew signal input
rlabel metal2 s 166814 359200 166870 359800 6 in[7]
port 108 nsew signal input
rlabel metal2 s 356150 359200 356206 359800 6 in[80]
port 109 nsew signal input
rlabel metal3 s 359200 118328 359800 118448 6 in[81]
port 110 nsew signal input
rlabel metal2 s 159730 200 159786 800 6 in[82]
port 111 nsew signal input
rlabel metal3 s 200 99288 800 99408 6 in[83]
port 112 nsew signal input
rlabel metal2 s 228638 200 228694 800 6 in[84]
port 113 nsew signal input
rlabel metal2 s 213826 200 213882 800 6 in[85]
port 114 nsew signal input
rlabel metal2 s 90822 200 90878 800 6 in[86]
port 115 nsew signal input
rlabel metal3 s 200 272008 800 272128 6 in[87]
port 116 nsew signal input
rlabel metal2 s 68926 200 68982 800 6 in[88]
port 117 nsew signal input
rlabel metal2 s 43810 359200 43866 359800 6 in[89]
port 118 nsew signal input
rlabel metal2 s 104990 200 105046 800 6 in[8]
port 119 nsew signal input
rlabel metal2 s 144918 200 144974 800 6 in[90]
port 120 nsew signal input
rlabel metal2 s 115938 200 115994 800 6 in[91]
port 121 nsew signal input
rlabel metal2 s 50250 200 50306 800 6 in[92]
port 122 nsew signal input
rlabel metal2 s 308494 200 308550 800 6 in[93]
port 123 nsew signal input
rlabel metal2 s 97906 200 97962 800 6 in[94]
port 124 nsew signal input
rlabel metal2 s 7102 359200 7158 359800 6 in[95]
port 125 nsew signal input
rlabel metal3 s 200 260448 800 260568 6 in[96]
port 126 nsew signal input
rlabel metal2 s 112718 359200 112774 359800 6 in[97]
port 127 nsew signal input
rlabel metal3 s 200 118328 800 118448 6 in[98]
port 128 nsew signal input
rlabel metal3 s 359200 348848 359800 348968 6 in[99]
port 129 nsew signal input
rlabel metal3 s 359200 133968 359800 134088 6 in[9]
port 130 nsew signal input
rlabel metal2 s 141698 200 141754 800 6 key[0]
port 131 nsew signal input
rlabel metal3 s 359200 53048 359800 53168 6 key[100]
port 132 nsew signal input
rlabel metal3 s 200 229848 800 229968 6 key[101]
port 133 nsew signal input
rlabel metal3 s 359200 38088 359800 38208 6 key[102]
port 134 nsew signal input
rlabel metal3 s 200 106768 800 106888 6 key[103]
port 135 nsew signal input
rlabel metal3 s 200 42168 800 42288 6 key[104]
port 136 nsew signal input
rlabel metal2 s 319442 200 319498 800 6 key[105]
port 137 nsew signal input
rlabel metal2 s 112074 200 112130 800 6 key[106]
port 138 nsew signal input
rlabel metal3 s 200 7488 800 7608 6 key[107]
port 139 nsew signal input
rlabel metal3 s 200 225768 800 225888 6 key[108]
port 140 nsew signal input
rlabel metal2 s 36082 359200 36138 359800 6 key[109]
port 141 nsew signal input
rlabel metal2 s 162950 200 163006 800 6 key[10]
port 142 nsew signal input
rlabel metal3 s 200 348848 800 348968 6 key[110]
port 143 nsew signal input
rlabel metal2 s 203522 359200 203578 359800 6 key[111]
port 144 nsew signal input
rlabel metal2 s 221554 359200 221610 359800 6 key[112]
port 145 nsew signal input
rlabel metal3 s 359200 321648 359800 321768 6 key[113]
port 146 nsew signal input
rlabel metal2 s 10966 359200 11022 359800 6 key[114]
port 147 nsew signal input
rlabel metal2 s 312358 359200 312414 359800 6 key[115]
port 148 nsew signal input
rlabel metal3 s 359200 122408 359800 122528 6 key[116]
port 149 nsew signal input
rlabel metal3 s 359200 129888 359800 130008 6 key[117]
port 150 nsew signal input
rlabel metal2 s 224774 200 224830 800 6 key[118]
port 151 nsew signal input
rlabel metal2 s 101126 200 101182 800 6 key[119]
port 152 nsew signal input
rlabel metal2 s 119802 200 119858 800 6 key[11]
port 153 nsew signal input
rlabel metal3 s 200 61208 800 61328 6 key[120]
port 154 nsew signal input
rlabel metal3 s 200 129888 800 130008 6 key[121]
port 155 nsew signal input
rlabel metal3 s 200 157088 800 157208 6 key[122]
port 156 nsew signal input
rlabel metal3 s 200 168648 800 168768 6 key[123]
port 157 nsew signal input
rlabel metal3 s 359200 233248 359800 233368 6 key[124]
port 158 nsew signal input
rlabel metal3 s 200 76168 800 76288 6 key[125]
port 159 nsew signal input
rlabel metal3 s 200 53048 800 53168 6 key[126]
port 160 nsew signal input
rlabel metal2 s 25134 359200 25190 359800 6 key[127]
port 161 nsew signal input
rlabel metal3 s 200 257048 800 257168 6 key[12]
port 162 nsew signal input
rlabel metal2 s 283378 359200 283434 359800 6 key[13]
port 163 nsew signal input
rlabel metal3 s 200 26528 800 26648 6 key[14]
port 164 nsew signal input
rlabel metal3 s 359200 57128 359800 57248 6 key[15]
port 165 nsew signal input
rlabel metal2 s 177762 359200 177818 359800 6 key[16]
port 166 nsew signal input
rlabel metal3 s 200 352928 800 353048 6 key[17]
port 167 nsew signal input
rlabel metal2 s 83738 359200 83794 359800 6 key[18]
port 168 nsew signal input
rlabel metal3 s 359200 229848 359800 229968 6 key[19]
port 169 nsew signal input
rlabel metal2 s 137834 200 137890 800 6 key[1]
port 170 nsew signal input
rlabel metal2 s 123022 200 123078 800 6 key[20]
port 171 nsew signal input
rlabel metal3 s 359200 114248 359800 114368 6 key[21]
port 172 nsew signal input
rlabel metal2 s 337474 200 337530 800 6 key[22]
port 173 nsew signal input
rlabel metal2 s 181626 359200 181682 359800 6 key[23]
port 174 nsew signal input
rlabel metal3 s 359200 22448 359800 22568 6 key[24]
port 175 nsew signal input
rlabel metal2 s 155866 200 155922 800 6 key[25]
port 176 nsew signal input
rlabel metal2 s 316222 359200 316278 359800 6 key[26]
port 177 nsew signal input
rlabel metal3 s 359200 237328 359800 237448 6 key[27]
port 178 nsew signal input
rlabel metal2 s 18 359200 74 359800 6 key[28]
port 179 nsew signal input
rlabel metal3 s 200 356328 800 356448 6 key[29]
port 180 nsew signal input
rlabel metal2 s 359370 359200 359426 359800 6 key[2]
port 181 nsew signal input
rlabel metal2 s 298190 359200 298246 359800 6 key[30]
port 182 nsew signal input
rlabel metal2 s 312358 200 312414 800 6 key[31]
port 183 nsew signal input
rlabel metal2 s 305274 359200 305330 359800 6 key[32]
port 184 nsew signal input
rlabel metal3 s 359200 252968 359800 253088 6 key[33]
port 185 nsew signal input
rlabel metal2 s 18050 200 18106 800 6 key[34]
port 186 nsew signal input
rlabel metal3 s 200 310768 800 310888 6 key[35]
port 187 nsew signal input
rlabel metal3 s 200 248888 800 249008 6 key[36]
port 188 nsew signal input
rlabel metal2 s 301410 200 301466 800 6 key[37]
port 189 nsew signal input
rlabel metal3 s 200 283568 800 283688 6 key[38]
port 190 nsew signal input
rlabel metal2 s 32862 359200 32918 359800 6 key[39]
port 191 nsew signal input
rlabel metal2 s 228638 359200 228694 359800 6 key[3]
port 192 nsew signal input
rlabel metal3 s 200 160488 800 160608 6 key[40]
port 193 nsew signal input
rlabel metal3 s 200 149608 800 149728 6 key[41]
port 194 nsew signal input
rlabel metal3 s 200 10888 800 11008 6 key[42]
port 195 nsew signal input
rlabel metal2 s 163594 359200 163650 359800 6 key[43]
port 196 nsew signal input
rlabel metal2 s 181626 200 181682 800 6 key[44]
port 197 nsew signal input
rlabel metal3 s 359200 202648 359800 202768 6 key[45]
port 198 nsew signal input
rlabel metal2 s 166814 200 166870 800 6 key[46]
port 199 nsew signal input
rlabel metal3 s 359200 48968 359800 49088 6 key[47]
port 200 nsew signal input
rlabel metal2 s 323306 359200 323362 359800 6 key[48]
port 201 nsew signal input
rlabel metal3 s 200 72768 800 72888 6 key[49]
port 202 nsew signal input
rlabel metal2 s 207386 359200 207442 359800 6 key[4]
port 203 nsew signal input
rlabel metal2 s 276294 359200 276350 359800 6 key[50]
port 204 nsew signal input
rlabel metal2 s 338118 359200 338174 359800 6 key[51]
port 205 nsew signal input
rlabel metal2 s 68926 359200 68982 359800 6 key[52]
port 206 nsew signal input
rlabel metal2 s 286598 200 286654 800 6 key[53]
port 207 nsew signal input
rlabel metal2 s 355506 200 355562 800 6 key[54]
port 208 nsew signal input
rlabel metal3 s 359200 68688 359800 68808 6 key[55]
port 209 nsew signal input
rlabel metal3 s 200 314168 800 314288 6 key[56]
port 210 nsew signal input
rlabel metal2 s 206742 200 206798 800 6 key[57]
port 211 nsew signal input
rlabel metal3 s 200 264528 800 264648 6 key[58]
port 212 nsew signal input
rlabel metal3 s 359200 99288 359800 99408 6 key[59]
port 213 nsew signal input
rlabel metal2 s 130750 359200 130806 359800 6 key[5]
port 214 nsew signal input
rlabel metal3 s 359200 167968 359800 168088 6 key[60]
port 215 nsew signal input
rlabel metal2 s 61842 359200 61898 359800 6 key[61]
port 216 nsew signal input
rlabel metal3 s 200 57128 800 57248 6 key[62]
port 217 nsew signal input
rlabel metal2 s 243450 200 243506 800 6 key[63]
port 218 nsew signal input
rlabel metal2 s 294326 200 294382 800 6 key[64]
port 219 nsew signal input
rlabel metal2 s 47030 200 47086 800 6 key[65]
port 220 nsew signal input
rlabel metal3 s 200 49648 800 49768 6 key[66]
port 221 nsew signal input
rlabel metal2 s 264702 200 264758 800 6 key[67]
port 222 nsew signal input
rlabel metal3 s 359200 3408 359800 3528 6 key[68]
port 223 nsew signal input
rlabel metal3 s 359200 153008 359800 153128 6 key[69]
port 224 nsew signal input
rlabel metal3 s 359200 352248 359800 352368 6 key[6]
port 225 nsew signal input
rlabel metal2 s 192574 359200 192630 359800 6 key[70]
port 226 nsew signal input
rlabel metal3 s 200 199248 800 199368 6 key[71]
port 227 nsew signal input
rlabel metal2 s 94042 200 94098 800 6 key[72]
port 228 nsew signal input
rlabel metal3 s 359200 191088 359800 191208 6 key[73]
port 229 nsew signal input
rlabel metal2 s 297546 200 297602 800 6 key[74]
port 230 nsew signal input
rlabel metal2 s 287242 359200 287298 359800 6 key[75]
port 231 nsew signal input
rlabel metal2 s 61198 200 61254 800 6 key[76]
port 232 nsew signal input
rlabel metal3 s 200 91808 800 91928 6 key[77]
port 233 nsew signal input
rlabel metal3 s 359200 310088 359800 310208 6 key[78]
port 234 nsew signal input
rlabel metal3 s 359200 329128 359800 329248 6 key[79]
port 235 nsew signal input
rlabel metal3 s 359200 279488 359800 279608 6 key[7]
port 236 nsew signal input
rlabel metal2 s 199658 359200 199714 359800 6 key[80]
port 237 nsew signal input
rlabel metal3 s 200 38088 800 38208 6 key[81]
port 238 nsew signal input
rlabel metal3 s 200 164568 800 164688 6 key[82]
port 239 nsew signal input
rlabel metal3 s 200 218288 800 218408 6 key[83]
port 240 nsew signal input
rlabel metal2 s 159730 359200 159786 359800 6 key[84]
port 241 nsew signal input
rlabel metal2 s 3238 200 3294 800 6 key[85]
port 242 nsew signal input
rlabel metal3 s 200 195168 800 195288 6 key[86]
port 243 nsew signal input
rlabel metal2 s 173898 200 173954 800 6 key[87]
port 244 nsew signal input
rlabel metal2 s 348422 200 348478 800 6 key[88]
port 245 nsew signal input
rlabel metal3 s 359200 344768 359800 344888 6 key[89]
port 246 nsew signal input
rlabel metal3 s 359200 18368 359800 18488 6 key[8]
port 247 nsew signal input
rlabel metal2 s 174542 359200 174598 359800 6 key[90]
port 248 nsew signal input
rlabel metal2 s 10322 200 10378 800 6 key[91]
port 249 nsew signal input
rlabel metal2 s 65062 200 65118 800 6 key[92]
port 250 nsew signal input
rlabel metal2 s 148782 200 148838 800 6 key[93]
port 251 nsew signal input
rlabel metal2 s 327170 359200 327226 359800 6 key[94]
port 252 nsew signal input
rlabel metal3 s 200 299208 800 299328 6 key[95]
port 253 nsew signal input
rlabel metal2 s 126886 200 126942 800 6 key[96]
port 254 nsew signal input
rlabel metal3 s 200 14968 800 15088 6 key[97]
port 255 nsew signal input
rlabel metal3 s 359200 148928 359800 149048 6 key[98]
port 256 nsew signal input
rlabel metal3 s 359200 218288 359800 218408 6 key[99]
port 257 nsew signal input
rlabel metal2 s 261482 200 261538 800 6 key[9]
port 258 nsew signal input
rlabel metal3 s 200 19048 800 19168 6 out[0]
port 259 nsew signal output
rlabel metal2 s 334254 200 334310 800 6 out[100]
port 260 nsew signal output
rlabel metal3 s 200 222368 800 222488 6 out[101]
port 261 nsew signal output
rlabel metal2 s 272430 359200 272486 359800 6 out[102]
port 262 nsew signal output
rlabel metal2 s 79874 359200 79930 359800 6 out[103]
port 263 nsew signal output
rlabel metal3 s 200 291048 800 291168 6 out[104]
port 264 nsew signal output
rlabel metal3 s 200 214208 800 214328 6 out[105]
port 265 nsew signal output
rlabel metal3 s 359200 14968 359800 15088 6 out[106]
port 266 nsew signal output
rlabel metal2 s 243450 359200 243506 359800 6 out[107]
port 267 nsew signal output
rlabel metal2 s 315578 200 315634 800 6 out[108]
port 268 nsew signal output
rlabel metal2 s 50894 359200 50950 359800 6 out[109]
port 269 nsew signal output
rlabel metal2 s 43166 200 43222 800 6 out[10]
port 270 nsew signal output
rlabel metal3 s 359200 160488 359800 160608 6 out[110]
port 271 nsew signal output
rlabel metal2 s 18050 359200 18106 359800 6 out[111]
port 272 nsew signal output
rlabel metal3 s 359200 214208 359800 214328 6 out[112]
port 273 nsew signal output
rlabel metal2 s 86958 200 87014 800 6 out[113]
port 274 nsew signal output
rlabel metal2 s 323306 200 323362 800 6 out[114]
port 275 nsew signal output
rlabel metal2 s 137834 359200 137890 359800 6 out[115]
port 276 nsew signal output
rlabel metal2 s 330390 359200 330446 359800 6 out[116]
port 277 nsew signal output
rlabel metal3 s 359200 256368 359800 256488 6 out[117]
port 278 nsew signal output
rlabel metal2 s 123666 359200 123722 359800 6 out[118]
port 279 nsew signal output
rlabel metal2 s 152646 359200 152702 359800 6 out[119]
port 280 nsew signal output
rlabel metal3 s 359200 45568 359800 45688 6 out[11]
port 281 nsew signal output
rlabel metal2 s 101770 359200 101826 359800 6 out[120]
port 282 nsew signal output
rlabel metal3 s 200 176128 800 176248 6 out[121]
port 283 nsew signal output
rlabel metal2 s 261482 359200 261538 359800 6 out[122]
port 284 nsew signal output
rlabel metal2 s 188710 359200 188766 359800 6 out[123]
port 285 nsew signal output
rlabel metal2 s 54758 359200 54814 359800 6 out[124]
port 286 nsew signal output
rlabel metal3 s 200 145528 800 145648 6 out[125]
port 287 nsew signal output
rlabel metal2 s 192574 200 192630 800 6 out[126]
port 288 nsew signal output
rlabel metal3 s 359200 248888 359800 249008 6 out[127]
port 289 nsew signal output
rlabel metal3 s 359200 225768 359800 225888 6 out[12]
port 290 nsew signal output
rlabel metal2 s 217690 200 217746 800 6 out[13]
port 291 nsew signal output
rlabel metal3 s 200 141448 800 141568 6 out[14]
port 292 nsew signal output
rlabel metal3 s 200 180208 800 180328 6 out[15]
port 293 nsew signal output
rlabel metal2 s 330390 200 330446 800 6 out[16]
port 294 nsew signal output
rlabel metal3 s 200 64608 800 64728 6 out[17]
port 295 nsew signal output
rlabel metal2 s 349066 359200 349122 359800 6 out[18]
port 296 nsew signal output
rlabel metal2 s 195794 200 195850 800 6 out[19]
port 297 nsew signal output
rlabel metal2 s 279514 200 279570 800 6 out[1]
port 298 nsew signal output
rlabel metal3 s 359200 64608 359800 64728 6 out[20]
port 299 nsew signal output
rlabel metal2 s 72790 359200 72846 359800 6 out[21]
port 300 nsew signal output
rlabel metal3 s 200 68688 800 68808 6 out[22]
port 301 nsew signal output
rlabel metal2 s 36082 200 36138 800 6 out[23]
port 302 nsew signal output
rlabel metal2 s 145562 359200 145618 359800 6 out[24]
port 303 nsew signal output
rlabel metal3 s 359200 195168 359800 195288 6 out[25]
port 304 nsew signal output
rlabel metal3 s 359200 333208 359800 333328 6 out[26]
port 305 nsew signal output
rlabel metal3 s 200 45568 800 45688 6 out[27]
port 306 nsew signal output
rlabel metal2 s 301410 359200 301466 359800 6 out[28]
port 307 nsew signal output
rlabel metal3 s 359200 137368 359800 137488 6 out[29]
port 308 nsew signal output
rlabel metal2 s 268566 200 268622 800 6 out[2]
port 309 nsew signal output
rlabel metal2 s 290462 359200 290518 359800 6 out[30]
port 310 nsew signal output
rlabel metal2 s 257618 200 257674 800 6 out[31]
port 311 nsew signal output
rlabel metal3 s 200 191768 800 191888 6 out[32]
port 312 nsew signal output
rlabel metal3 s 200 252968 800 253088 6 out[33]
port 313 nsew signal output
rlabel metal2 s 345202 200 345258 800 6 out[34]
port 314 nsew signal output
rlabel metal3 s 359200 83648 359800 83768 6 out[35]
port 315 nsew signal output
rlabel metal2 s 134614 359200 134670 359800 6 out[36]
port 316 nsew signal output
rlabel metal3 s 359200 302608 359800 302728 6 out[37]
port 317 nsew signal output
rlabel metal3 s 200 302608 800 302728 6 out[38]
port 318 nsew signal output
rlabel metal3 s 200 329808 800 329928 6 out[39]
port 319 nsew signal output
rlabel metal3 s 200 318248 800 318368 6 out[3]
port 320 nsew signal output
rlabel metal2 s 14186 200 14242 800 6 out[40]
port 321 nsew signal output
rlabel metal3 s 200 84328 800 84448 6 out[41]
port 322 nsew signal output
rlabel metal3 s 359200 176128 359800 176248 6 out[42]
port 323 nsew signal output
rlabel metal2 s 199658 200 199714 800 6 out[43]
port 324 nsew signal output
rlabel metal2 s 258262 359200 258318 359800 6 out[44]
port 325 nsew signal output
rlabel metal2 s 341338 359200 341394 359800 6 out[45]
port 326 nsew signal output
rlabel metal2 s 39946 359200 40002 359800 6 out[46]
port 327 nsew signal output
rlabel metal2 s 54114 200 54170 800 6 out[47]
port 328 nsew signal output
rlabel metal3 s 359200 206728 359800 206848 6 out[48]
port 329 nsew signal output
rlabel metal2 s 352286 359200 352342 359800 6 out[49]
port 330 nsew signal output
rlabel metal3 s 200 233928 800 234048 6 out[4]
port 331 nsew signal output
rlabel metal3 s 359200 272008 359800 272128 6 out[50]
port 332 nsew signal output
rlabel metal3 s 359200 106768 359800 106888 6 out[51]
port 333 nsew signal output
rlabel metal2 s 239586 200 239642 800 6 out[52]
port 334 nsew signal output
rlabel metal2 s 309138 359200 309194 359800 6 out[53]
port 335 nsew signal output
rlabel metal2 s 105634 359200 105690 359800 6 out[54]
port 336 nsew signal output
rlabel metal2 s 108854 200 108910 800 6 out[55]
port 337 nsew signal output
rlabel metal3 s 359200 210128 359800 210248 6 out[56]
port 338 nsew signal output
rlabel metal2 s 283378 200 283434 800 6 out[57]
port 339 nsew signal output
rlabel metal3 s 359200 95208 359800 95328 6 out[58]
port 340 nsew signal output
rlabel metal3 s 200 206728 800 206848 6 out[59]
port 341 nsew signal output
rlabel metal2 s 359370 200 359426 800 6 out[5]
port 342 nsew signal output
rlabel metal2 s 57978 200 58034 800 6 out[60]
port 343 nsew signal output
rlabel metal2 s 170678 200 170734 800 6 out[61]
port 344 nsew signal output
rlabel metal3 s 359200 145528 359800 145648 6 out[62]
port 345 nsew signal output
rlabel metal2 s 294326 359200 294382 359800 6 out[63]
port 346 nsew signal output
rlabel metal3 s 359200 317568 359800 317688 6 out[64]
port 347 nsew signal output
rlabel metal3 s 359200 6808 359800 6928 6 out[65]
port 348 nsew signal output
rlabel metal2 s 28998 200 29054 800 6 out[66]
port 349 nsew signal output
rlabel metal3 s 359200 199248 359800 199368 6 out[67]
port 350 nsew signal output
rlabel metal2 s 7102 200 7158 800 6 out[68]
port 351 nsew signal output
rlabel metal3 s 359200 325728 359800 325848 6 out[69]
port 352 nsew signal output
rlabel metal2 s 279514 359200 279570 359800 6 out[6]
port 353 nsew signal output
rlabel metal3 s 359200 29928 359800 30048 6 out[70]
port 354 nsew signal output
rlabel metal2 s 265346 359200 265402 359800 6 out[71]
port 355 nsew signal output
rlabel metal3 s 200 110848 800 110968 6 out[72]
port 356 nsew signal output
rlabel metal3 s 200 122408 800 122528 6 out[73]
port 357 nsew signal output
rlabel metal2 s 235722 200 235778 800 6 out[74]
port 358 nsew signal output
rlabel metal2 s 18 200 74 800 6 out[75]
port 359 nsew signal output
rlabel metal2 s 275650 200 275706 800 6 out[76]
port 360 nsew signal output
rlabel metal3 s 200 183608 800 183728 6 out[77]
port 361 nsew signal output
rlabel metal3 s 200 325728 800 325848 6 out[78]
port 362 nsew signal output
rlabel metal2 s 108854 359200 108910 359800 6 out[79]
port 363 nsew signal output
rlabel metal3 s 200 126488 800 126608 6 out[7]
port 364 nsew signal output
rlabel metal2 s 72146 200 72202 800 6 out[80]
port 365 nsew signal output
rlabel metal2 s 25134 200 25190 800 6 out[81]
port 366 nsew signal output
rlabel metal2 s 196438 359200 196494 359800 6 out[82]
port 367 nsew signal output
rlabel metal2 s 115938 359200 115994 359800 6 out[83]
port 368 nsew signal output
rlabel metal2 s 188710 200 188766 800 6 out[84]
port 369 nsew signal output
rlabel metal2 s 254398 359200 254454 359800 6 out[85]
port 370 nsew signal output
rlabel metal3 s 359200 91808 359800 91928 6 out[86]
port 371 nsew signal output
rlabel metal3 s 200 245488 800 245608 6 out[87]
port 372 nsew signal output
rlabel metal3 s 359200 275408 359800 275528 6 out[88]
port 373 nsew signal output
rlabel metal2 s 76010 200 76066 800 6 out[89]
port 374 nsew signal output
rlabel metal2 s 133970 200 134026 800 6 out[8]
port 375 nsew signal output
rlabel metal3 s 200 34008 800 34128 6 out[90]
port 376 nsew signal output
rlabel metal3 s 359200 263848 359800 263968 6 out[91]
port 377 nsew signal output
rlabel metal2 s 210606 200 210662 800 6 out[92]
port 378 nsew signal output
rlabel metal2 s 239586 359200 239642 359800 6 out[93]
port 379 nsew signal output
rlabel metal2 s 236366 359200 236422 359800 6 out[94]
port 380 nsew signal output
rlabel metal3 s 200 341368 800 341488 6 out[95]
port 381 nsew signal output
rlabel metal2 s 47030 359200 47086 359800 6 out[96]
port 382 nsew signal output
rlabel metal2 s 253754 200 253810 800 6 out[97]
port 383 nsew signal output
rlabel metal3 s 200 80248 800 80368 6 out[98]
port 384 nsew signal output
rlabel metal3 s 200 306688 800 306808 6 out[99]
port 385 nsew signal output
rlabel metal3 s 359200 172048 359800 172168 6 out[9]
port 386 nsew signal output
rlabel metal4 s 4208 2128 4528 357456 6 vccd1
port 387 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 357456 6 vccd1
port 387 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 357456 6 vccd1
port 387 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 357456 6 vccd1
port 387 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 357456 6 vccd1
port 387 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 357456 6 vccd1
port 387 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 357456 6 vccd1
port 387 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 357456 6 vccd1
port 387 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 357456 6 vccd1
port 387 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 357456 6 vccd1
port 387 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 357456 6 vccd1
port 387 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 357456 6 vccd1
port 387 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 357456 6 vssd1
port 388 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 357456 6 vssd1
port 388 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 357456 6 vssd1
port 388 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 357456 6 vssd1
port 388 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 357456 6 vssd1
port 388 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 357456 6 vssd1
port 388 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 357456 6 vssd1
port 388 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 357456 6 vssd1
port 388 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 357456 6 vssd1
port 388 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 357456 6 vssd1
port 388 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 357456 6 vssd1
port 388 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 357456 6 vssd1
port 388 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 360000 360000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 209165004
string GDS_FILE /home/urielcho/Proyectos_caravel/MPW8/decrypt_aes128/openlane/decrypt_aes128/runs/22_12_20_18_34/results/signoff/decrypt_aes128.magic.gds
string GDS_START 1459838
<< end >>

