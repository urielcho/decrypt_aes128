VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO decrypt_aes128
  CLASS BLOCK ;
  FOREIGN decrypt_aes128 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1800.000 BY 1800.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1492.640 1799.000 1493.240 ;
    END
  END clk
  PIN decReset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1706.690 1.000 1706.970 4.000 ;
    END
  END decReset
  PIN in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 170.040 1799.000 170.640 ;
    END
  END in[0]
  PIN in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1666.040 4.000 1666.640 ;
    END
  END in[100]
  PIN in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1686.440 4.000 1687.040 ;
    END
  END in[101]
  PIN in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1452.310 1.000 1452.590 4.000 ;
    END
  END in[102]
  PIN in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 360.440 1799.000 361.040 ;
    END
  END in[103]
  PIN in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 1796.000 927.730 1799.000 ;
    END
  END in[104]
  PIN in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 153.040 4.000 153.640 ;
    END
  END in[105]
  PIN in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1207.040 4.000 1207.640 ;
    END
  END in[106]
  PIN in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 1796.000 744.190 1799.000 ;
    END
  END in[107]
  PIN in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 1796.000 1072.630 1799.000 ;
    END
  END in[108]
  PIN in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1236.570 1796.000 1236.850 1799.000 ;
    END
  END in[109]
  PIN in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 1796.000 435.070 1799.000 ;
    END
  END in[10]
  PIN in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.210 1796.000 1597.490 1799.000 ;
    END
  END in[110]
  PIN in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 479.440 4.000 480.040 ;
    END
  END in[111]
  PIN in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1761.430 1.000 1761.710 4.000 ;
    END
  END in[112]
  PIN in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 1.000 399.650 4.000 ;
    END
  END in[113]
  PIN in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1054.040 4.000 1054.640 ;
    END
  END in[114]
  PIN in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1016.640 4.000 1017.240 ;
    END
  END in[115]
  PIN in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.830 1796.000 1343.110 1799.000 ;
    END
  END in[116]
  PIN in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1703.440 1799.000 1704.040 ;
    END
  END in[117]
  PIN in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 1796.000 325.590 1799.000 ;
    END
  END in[118]
  PIN in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 513.440 1799.000 514.040 ;
    END
  END in[119]
  PIN in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1475.640 4.000 1476.240 ;
    END
  END in[11]
  PIN in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1108.440 1799.000 1109.040 ;
    END
  END in[120]
  PIN in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.150 1.000 1362.430 4.000 ;
    END
  END in[121]
  PIN in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 1.000 654.030 4.000 ;
    END
  END in[122]
  PIN in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 1796.000 599.290 1799.000 ;
    END
  END in[123]
  PIN in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 897.640 1799.000 898.240 ;
    END
  END in[124]
  PIN in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.350 1.000 1233.630 4.000 ;
    END
  END in[125]
  PIN in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1302.240 1799.000 1302.840 ;
    END
  END in[126]
  PIN in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1339.640 1799.000 1340.240 ;
    END
  END in[127]
  PIN in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 1.000 415.750 4.000 ;
    END
  END in[12]
  PIN in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 938.440 1799.000 939.040 ;
    END
  END in[13]
  PIN in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 1.000 106.630 4.000 ;
    END
  END in[14]
  PIN in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1397.440 4.000 1398.040 ;
    END
  END in[15]
  PIN in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1339.640 4.000 1340.240 ;
    END
  END in[16]
  PIN in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 574.640 4.000 575.240 ;
    END
  END in[17]
  PIN in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1608.240 4.000 1608.840 ;
    END
  END in[18]
  PIN in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.010 1796.000 1726.290 1799.000 ;
    END
  END in[19]
  PIN in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 554.240 1799.000 554.840 ;
    END
  END in[1]
  PIN in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 1.000 1162.790 4.000 ;
    END
  END in[20]
  PIN in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1207.040 1799.000 1207.640 ;
    END
  END in[21]
  PIN in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.230 1.000 924.510 4.000 ;
    END
  END in[22]
  PIN in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1781.640 1799.000 1782.240 ;
    END
  END in[23]
  PIN in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.670 1796.000 1252.950 1799.000 ;
    END
  END in[24]
  PIN in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 1796.000 19.690 1799.000 ;
    END
  END in[25]
  PIN in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 112.240 4.000 112.840 ;
    END
  END in[26]
  PIN in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 707.240 1799.000 707.840 ;
    END
  END in[27]
  PIN in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 438.640 1799.000 439.240 ;
    END
  END in[28]
  PIN in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 1.000 161.370 4.000 ;
    END
  END in[29]
  PIN in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 938.440 4.000 939.040 ;
    END
  END in[2]
  PIN in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 17.040 4.000 17.640 ;
    END
  END in[30]
  PIN in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 1796.000 109.850 1799.000 ;
    END
  END in[31]
  PIN in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1533.440 1799.000 1534.040 ;
    END
  END in[32]
  PIN in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.450 1796.000 1088.730 1799.000 ;
    END
  END in[33]
  PIN in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 1796.000 634.710 1799.000 ;
    END
  END in[34]
  PIN in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 669.840 4.000 670.440 ;
    END
  END in[35]
  PIN in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 401.240 1799.000 401.840 ;
    END
  END in[36]
  PIN in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 782.040 1799.000 782.640 ;
    END
  END in[37]
  PIN in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 918.040 1799.000 918.640 ;
    END
  END in[38]
  PIN in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.770 1.000 1108.050 4.000 ;
    END
  END in[39]
  PIN in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 380.840 1799.000 381.440 ;
    END
  END in[3]
  PIN in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 765.040 4.000 765.640 ;
    END
  END in[40]
  PIN in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 1796.000 454.390 1799.000 ;
    END
  END in[41]
  PIN in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.150 1.000 1523.430 4.000 ;
    END
  END in[42]
  PIN in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1186.640 4.000 1187.240 ;
    END
  END in[43]
  PIN in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.670 1.000 1252.950 4.000 ;
    END
  END in[44]
  PIN in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 1796.000 1127.370 1799.000 ;
    END
  END in[45]
  PIN in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 1796.000 489.810 1799.000 ;
    END
  END in[46]
  PIN in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1723.840 4.000 1724.440 ;
    END
  END in[47]
  PIN in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.030 1796.000 1053.310 1799.000 ;
    END
  END in[48]
  PIN in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 1.000 889.090 4.000 ;
    END
  END in[49]
  PIN in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 207.440 1799.000 208.040 ;
    END
  END in[4]
  PIN in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 1796.000 782.830 1799.000 ;
    END
  END in[50]
  PIN in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 1.000 760.290 4.000 ;
    END
  END in[51]
  PIN in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 516.840 4.000 517.440 ;
    END
  END in[52]
  PIN in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 1796.000 708.770 1799.000 ;
    END
  END in[53]
  PIN in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 1796.000 1162.790 1799.000 ;
    END
  END in[54]
  PIN in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1455.240 1799.000 1455.840 ;
    END
  END in[55]
  PIN in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 1.000 200.010 4.000 ;
    END
  END in[56]
  PIN in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.390 1.000 1014.670 4.000 ;
    END
  END in[57]
  PIN in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1686.440 1799.000 1687.040 ;
    END
  END in[58]
  PIN in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 1796.000 380.330 1799.000 ;
    END
  END in[59]
  PIN in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.270 1796.000 1671.550 1799.000 ;
    END
  END in[5]
  PIN in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 860.240 4.000 860.840 ;
    END
  END in[60]
  PIN in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1475.640 1799.000 1476.240 ;
    END
  END in[61]
  PIN in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 690.240 4.000 690.840 ;
    END
  END in[62]
  PIN in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 1796.000 853.670 1799.000 ;
    END
  END in[63]
  PIN in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 302.640 1799.000 303.240 ;
    END
  END in[64]
  PIN in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 629.040 1799.000 629.640 ;
    END
  END in[65]
  PIN in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.630 1.000 1632.910 4.000 ;
    END
  END in[66]
  PIN in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1570.840 1799.000 1571.440 ;
    END
  END in[67]
  PIN in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 438.640 4.000 439.240 ;
    END
  END in[68]
  PIN in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 1796.000 145.270 1799.000 ;
    END
  END in[69]
  PIN in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 1796.000 473.710 1799.000 ;
    END
  END in[6]
  PIN in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 132.640 1799.000 133.240 ;
    END
  END in[70]
  PIN in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1380.440 4.000 1381.040 ;
    END
  END in[71]
  PIN in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1438.240 4.000 1438.840 ;
    END
  END in[72]
  PIN in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1434.840 1799.000 1435.440 ;
    END
  END in[73]
  PIN in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 822.840 1799.000 823.440 ;
    END
  END in[74]
  PIN in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1417.840 1799.000 1418.440 ;
    END
  END in[75]
  PIN in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1224.040 1799.000 1224.640 ;
    END
  END in[76]
  PIN in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 1796.000 71.210 1799.000 ;
    END
  END in[77]
  PIN in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 54.440 1799.000 55.040 ;
    END
  END in[78]
  PIN in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 1796.000 290.170 1799.000 ;
    END
  END in[79]
  PIN in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 1796.000 834.350 1799.000 ;
    END
  END in[7]
  PIN in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1780.750 1796.000 1781.030 1799.000 ;
    END
  END in[80]
  PIN in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 591.640 1799.000 592.240 ;
    END
  END in[81]
  PIN in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 1.000 798.930 4.000 ;
    END
  END in[82]
  PIN in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 496.440 4.000 497.040 ;
    END
  END in[83]
  PIN in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.190 1.000 1143.470 4.000 ;
    END
  END in[84]
  PIN in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.130 1.000 1069.410 4.000 ;
    END
  END in[85]
  PIN in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 1.000 454.390 4.000 ;
    END
  END in[86]
  PIN in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1360.040 4.000 1360.640 ;
    END
  END in[87]
  PIN in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 1.000 344.910 4.000 ;
    END
  END in[88]
  PIN in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 1796.000 219.330 1799.000 ;
    END
  END in[89]
  PIN in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 1.000 525.230 4.000 ;
    END
  END in[8]
  PIN in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 1.000 724.870 4.000 ;
    END
  END in[90]
  PIN in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 1.000 579.970 4.000 ;
    END
  END in[91]
  PIN in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 1.000 251.530 4.000 ;
    END
  END in[92]
  PIN in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.470 1.000 1542.750 4.000 ;
    END
  END in[93]
  PIN in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 1.000 489.810 4.000 ;
    END
  END in[94]
  PIN in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 1796.000 35.790 1799.000 ;
    END
  END in[95]
  PIN in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1302.240 4.000 1302.840 ;
    END
  END in[96]
  PIN in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 1796.000 563.870 1799.000 ;
    END
  END in[97]
  PIN in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 591.640 4.000 592.240 ;
    END
  END in[98]
  PIN in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1744.240 1799.000 1744.840 ;
    END
  END in[99]
  PIN in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 669.840 1799.000 670.440 ;
    END
  END in[9]
  PIN key[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 1.000 708.770 4.000 ;
    END
  END key[0]
  PIN key[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 265.240 1799.000 265.840 ;
    END
  END key[100]
  PIN key[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1149.240 4.000 1149.840 ;
    END
  END key[101]
  PIN key[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 190.440 1799.000 191.040 ;
    END
  END key[102]
  PIN key[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 533.840 4.000 534.440 ;
    END
  END key[103]
  PIN key[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 210.840 4.000 211.440 ;
    END
  END key[104]
  PIN key[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.210 1.000 1597.490 4.000 ;
    END
  END key[105]
  PIN key[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 1.000 560.650 4.000 ;
    END
  END key[106]
  PIN key[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 37.440 4.000 38.040 ;
    END
  END key[107]
  PIN key[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1128.840 4.000 1129.440 ;
    END
  END key[108]
  PIN key[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 1796.000 180.690 1799.000 ;
    END
  END key[109]
  PIN key[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.750 1.000 815.030 4.000 ;
    END
  END key[10]
  PIN key[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1744.240 4.000 1744.840 ;
    END
  END key[110]
  PIN key[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.610 1796.000 1017.890 1799.000 ;
    END
  END key[111]
  PIN key[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.770 1796.000 1108.050 1799.000 ;
    END
  END key[112]
  PIN key[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1608.240 1799.000 1608.840 ;
    END
  END key[113]
  PIN key[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 1796.000 55.110 1799.000 ;
    END
  END key[114]
  PIN key[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.790 1796.000 1562.070 1799.000 ;
    END
  END key[115]
  PIN key[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 612.040 1799.000 612.640 ;
    END
  END key[116]
  PIN key[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 649.440 1799.000 650.040 ;
    END
  END key[117]
  PIN key[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.870 1.000 1124.150 4.000 ;
    END
  END key[118]
  PIN key[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 1.000 505.910 4.000 ;
    END
  END key[119]
  PIN key[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 1.000 599.290 4.000 ;
    END
  END key[11]
  PIN key[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 306.040 4.000 306.640 ;
    END
  END key[120]
  PIN key[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 649.440 4.000 650.040 ;
    END
  END key[121]
  PIN key[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 785.440 4.000 786.040 ;
    END
  END key[122]
  PIN key[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 843.240 4.000 843.840 ;
    END
  END key[123]
  PIN key[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1166.240 1799.000 1166.840 ;
    END
  END key[124]
  PIN key[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 380.840 4.000 381.440 ;
    END
  END key[125]
  PIN key[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 265.240 4.000 265.840 ;
    END
  END key[126]
  PIN key[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 1796.000 125.950 1799.000 ;
    END
  END key[127]
  PIN key[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1285.240 4.000 1285.840 ;
    END
  END key[12]
  PIN key[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.890 1796.000 1417.170 1799.000 ;
    END
  END key[13]
  PIN key[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 132.640 4.000 133.240 ;
    END
  END key[14]
  PIN key[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 285.640 1799.000 286.240 ;
    END
  END key[15]
  PIN key[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 1796.000 889.090 1799.000 ;
    END
  END key[16]
  PIN key[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1764.640 4.000 1765.240 ;
    END
  END key[17]
  PIN key[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 1796.000 418.970 1799.000 ;
    END
  END key[18]
  PIN key[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1149.240 1799.000 1149.840 ;
    END
  END key[19]
  PIN key[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 1.000 689.450 4.000 ;
    END
  END key[1]
  PIN key[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 1.000 615.390 4.000 ;
    END
  END key[20]
  PIN key[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 571.240 1799.000 571.840 ;
    END
  END key[21]
  PIN key[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.370 1.000 1687.650 4.000 ;
    END
  END key[22]
  PIN key[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130 1796.000 908.410 1799.000 ;
    END
  END key[23]
  PIN key[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 112.240 1799.000 112.840 ;
    END
  END key[24]
  PIN key[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 1.000 779.610 4.000 ;
    END
  END key[25]
  PIN key[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.110 1796.000 1581.390 1799.000 ;
    END
  END key[26]
  PIN key[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1186.640 1799.000 1187.240 ;
    END
  END key[27]
  PIN key[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 1796.000 0.370 1799.000 ;
    END
  END key[28]
  PIN key[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1781.640 4.000 1782.240 ;
    END
  END key[29]
  PIN key[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1796.850 1796.000 1797.130 1799.000 ;
    END
  END key[2]
  PIN key[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 1796.000 1491.230 1799.000 ;
    END
  END key[30]
  PIN key[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.790 1.000 1562.070 4.000 ;
    END
  END key[31]
  PIN key[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.370 1796.000 1526.650 1799.000 ;
    END
  END key[32]
  PIN key[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1264.840 1799.000 1265.440 ;
    END
  END key[33]
  PIN key[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 1.000 90.530 4.000 ;
    END
  END key[34]
  PIN key[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1553.840 4.000 1554.440 ;
    END
  END key[35]
  PIN key[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1244.440 4.000 1245.040 ;
    END
  END key[36]
  PIN key[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.050 1.000 1507.330 4.000 ;
    END
  END key[37]
  PIN key[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1417.840 4.000 1418.440 ;
    END
  END key[38]
  PIN key[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 1796.000 164.590 1799.000 ;
    END
  END key[39]
  PIN key[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.190 1796.000 1143.470 1799.000 ;
    END
  END key[3]
  PIN key[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 802.440 4.000 803.040 ;
    END
  END key[40]
  PIN key[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 748.040 4.000 748.640 ;
    END
  END key[41]
  PIN key[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 54.440 4.000 55.040 ;
    END
  END key[42]
  PIN key[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 1796.000 818.250 1799.000 ;
    END
  END key[43]
  PIN key[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130 1.000 908.410 4.000 ;
    END
  END key[44]
  PIN key[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1013.240 1799.000 1013.840 ;
    END
  END key[45]
  PIN key[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 1.000 834.350 4.000 ;
    END
  END key[46]
  PIN key[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 244.840 1799.000 245.440 ;
    END
  END key[47]
  PIN key[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.530 1796.000 1616.810 1799.000 ;
    END
  END key[48]
  PIN key[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 363.840 4.000 364.440 ;
    END
  END key[49]
  PIN key[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.930 1796.000 1037.210 1799.000 ;
    END
  END key[4]
  PIN key[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.470 1796.000 1381.750 1799.000 ;
    END
  END key[50]
  PIN key[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1690.590 1796.000 1690.870 1799.000 ;
    END
  END key[51]
  PIN key[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 1796.000 344.910 1799.000 ;
    END
  END key[52]
  PIN key[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.990 1.000 1433.270 4.000 ;
    END
  END key[53]
  PIN key[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.530 1.000 1777.810 4.000 ;
    END
  END key[54]
  PIN key[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 343.440 1799.000 344.040 ;
    END
  END key[55]
  PIN key[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1570.840 4.000 1571.440 ;
    END
  END key[56]
  PIN key[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 1.000 1033.990 4.000 ;
    END
  END key[57]
  PIN key[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1322.640 4.000 1323.240 ;
    END
  END key[58]
  PIN key[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 496.440 1799.000 497.040 ;
    END
  END key[59]
  PIN key[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 1796.000 654.030 1799.000 ;
    END
  END key[5]
  PIN key[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 839.840 1799.000 840.440 ;
    END
  END key[60]
  PIN key[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 1796.000 309.490 1799.000 ;
    END
  END key[61]
  PIN key[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 285.640 4.000 286.240 ;
    END
  END key[62]
  PIN key[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.250 1.000 1217.530 4.000 ;
    END
  END key[63]
  PIN key[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.630 1.000 1471.910 4.000 ;
    END
  END key[64]
  PIN key[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 1.000 235.430 4.000 ;
    END
  END key[65]
  PIN key[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 248.240 4.000 248.840 ;
    END
  END key[66]
  PIN key[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.510 1.000 1323.790 4.000 ;
    END
  END key[67]
  PIN key[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 17.040 1799.000 17.640 ;
    END
  END key[68]
  PIN key[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 765.040 1799.000 765.640 ;
    END
  END key[69]
  PIN key[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1761.240 1799.000 1761.840 ;
    END
  END key[6]
  PIN key[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 1796.000 963.150 1799.000 ;
    END
  END key[70]
  PIN key[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 996.240 4.000 996.840 ;
    END
  END key[71]
  PIN key[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 1.000 470.490 4.000 ;
    END
  END key[72]
  PIN key[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 955.440 1799.000 956.040 ;
    END
  END key[73]
  PIN key[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1487.730 1.000 1488.010 4.000 ;
    END
  END key[74]
  PIN key[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.210 1796.000 1436.490 1799.000 ;
    END
  END key[75]
  PIN key[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 1.000 306.270 4.000 ;
    END
  END key[76]
  PIN key[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 459.040 4.000 459.640 ;
    END
  END key[77]
  PIN key[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1550.440 1799.000 1551.040 ;
    END
  END key[78]
  PIN key[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1645.640 1799.000 1646.240 ;
    END
  END key[79]
  PIN key[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1397.440 1799.000 1398.040 ;
    END
  END key[7]
  PIN key[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.290 1796.000 998.570 1799.000 ;
    END
  END key[80]
  PIN key[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 190.440 4.000 191.040 ;
    END
  END key[81]
  PIN key[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 822.840 4.000 823.440 ;
    END
  END key[82]
  PIN key[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1091.440 4.000 1092.040 ;
    END
  END key[83]
  PIN key[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 1796.000 798.930 1799.000 ;
    END
  END key[84]
  PIN key[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 1.000 16.470 4.000 ;
    END
  END key[85]
  PIN key[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 975.840 4.000 976.440 ;
    END
  END key[86]
  PIN key[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 1.000 869.770 4.000 ;
    END
  END key[87]
  PIN key[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.110 1.000 1742.390 4.000 ;
    END
  END key[88]
  PIN key[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1723.840 1799.000 1724.440 ;
    END
  END key[89]
  PIN key[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 91.840 1799.000 92.440 ;
    END
  END key[8]
  PIN key[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 1796.000 872.990 1799.000 ;
    END
  END key[90]
  PIN key[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 1.000 51.890 4.000 ;
    END
  END key[91]
  PIN key[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 1.000 325.590 4.000 ;
    END
  END key[92]
  PIN key[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 1.000 744.190 4.000 ;
    END
  END key[93]
  PIN key[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1635.850 1796.000 1636.130 1799.000 ;
    END
  END key[94]
  PIN key[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1496.040 4.000 1496.640 ;
    END
  END key[95]
  PIN key[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 1.000 634.710 4.000 ;
    END
  END key[96]
  PIN key[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 74.840 4.000 75.440 ;
    END
  END key[97]
  PIN key[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 744.640 1799.000 745.240 ;
    END
  END key[98]
  PIN key[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1091.440 1799.000 1092.040 ;
    END
  END key[99]
  PIN key[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.410 1.000 1307.690 4.000 ;
    END
  END key[9]
  PIN out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 95.240 4.000 95.840 ;
    END
  END out[0]
  PIN out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.270 1.000 1671.550 4.000 ;
    END
  END out[100]
  PIN out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1111.840 4.000 1112.440 ;
    END
  END out[101]
  PIN out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.150 1796.000 1362.430 1799.000 ;
    END
  END out[102]
  PIN out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 1796.000 399.650 1799.000 ;
    END
  END out[103]
  PIN out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1455.240 4.000 1455.840 ;
    END
  END out[104]
  PIN out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1071.040 4.000 1071.640 ;
    END
  END out[105]
  PIN out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 74.840 1799.000 75.440 ;
    END
  END out[106]
  PIN out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.250 1796.000 1217.530 1799.000 ;
    END
  END out[107]
  PIN out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1577.890 1.000 1578.170 4.000 ;
    END
  END out[108]
  PIN out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 1796.000 254.750 1799.000 ;
    END
  END out[109]
  PIN out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 1.000 216.110 4.000 ;
    END
  END out[10]
  PIN out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 802.440 1799.000 803.040 ;
    END
  END out[110]
  PIN out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 1796.000 90.530 1799.000 ;
    END
  END out[111]
  PIN out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1071.040 1799.000 1071.640 ;
    END
  END out[112]
  PIN out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 1.000 435.070 4.000 ;
    END
  END out[113]
  PIN out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.530 1.000 1616.810 4.000 ;
    END
  END out[114]
  PIN out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 1796.000 689.450 1799.000 ;
    END
  END out[115]
  PIN out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.950 1796.000 1652.230 1799.000 ;
    END
  END out[116]
  PIN out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1281.840 1799.000 1282.440 ;
    END
  END out[117]
  PIN out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 1796.000 618.610 1799.000 ;
    END
  END out[118]
  PIN out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 1796.000 763.510 1799.000 ;
    END
  END out[119]
  PIN out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 227.840 1799.000 228.440 ;
    END
  END out[11]
  PIN out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 1796.000 509.130 1799.000 ;
    END
  END out[120]
  PIN out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 880.640 4.000 881.240 ;
    END
  END out[121]
  PIN out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.410 1796.000 1307.690 1799.000 ;
    END
  END out[122]
  PIN out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 1796.000 943.830 1799.000 ;
    END
  END out[123]
  PIN out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 1796.000 274.070 1799.000 ;
    END
  END out[124]
  PIN out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 727.640 4.000 728.240 ;
    END
  END out[125]
  PIN out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 1.000 963.150 4.000 ;
    END
  END out[126]
  PIN out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1244.440 1799.000 1245.040 ;
    END
  END out[127]
  PIN out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1128.840 1799.000 1129.440 ;
    END
  END out[12]
  PIN out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.450 1.000 1088.730 4.000 ;
    END
  END out[13]
  PIN out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 707.240 4.000 707.840 ;
    END
  END out[14]
  PIN out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 901.040 4.000 901.640 ;
    END
  END out[15]
  PIN out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.950 1.000 1652.230 4.000 ;
    END
  END out[16]
  PIN out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 323.040 4.000 323.640 ;
    END
  END out[17]
  PIN out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.330 1796.000 1745.610 1799.000 ;
    END
  END out[18]
  PIN out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 1.000 979.250 4.000 ;
    END
  END out[19]
  PIN out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.570 1.000 1397.850 4.000 ;
    END
  END out[1]
  PIN out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 323.040 1799.000 323.640 ;
    END
  END out[20]
  PIN out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 1796.000 364.230 1799.000 ;
    END
  END out[21]
  PIN out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 343.440 4.000 344.040 ;
    END
  END out[22]
  PIN out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 1.000 180.690 4.000 ;
    END
  END out[23]
  PIN out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 1796.000 728.090 1799.000 ;
    END
  END out[24]
  PIN out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 975.840 1799.000 976.440 ;
    END
  END out[25]
  PIN out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1666.040 1799.000 1666.640 ;
    END
  END out[26]
  PIN out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 227.840 4.000 228.440 ;
    END
  END out[27]
  PIN out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.050 1796.000 1507.330 1799.000 ;
    END
  END out[28]
  PIN out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 686.840 1799.000 687.440 ;
    END
  END out[29]
  PIN out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.830 1.000 1343.110 4.000 ;
    END
  END out[2]
  PIN out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1452.310 1796.000 1452.590 1799.000 ;
    END
  END out[30]
  PIN out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1288.090 1.000 1288.370 4.000 ;
    END
  END out[31]
  PIN out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 958.840 4.000 959.440 ;
    END
  END out[32]
  PIN out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1264.840 4.000 1265.440 ;
    END
  END out[33]
  PIN out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.010 1.000 1726.290 4.000 ;
    END
  END out[34]
  PIN out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 418.240 1799.000 418.840 ;
    END
  END out[35]
  PIN out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 1796.000 673.350 1799.000 ;
    END
  END out[36]
  PIN out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1513.040 1799.000 1513.640 ;
    END
  END out[37]
  PIN out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1513.040 4.000 1513.640 ;
    END
  END out[38]
  PIN out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1649.040 4.000 1649.640 ;
    END
  END out[39]
  PIN out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1591.240 4.000 1591.840 ;
    END
  END out[3]
  PIN out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 1.000 71.210 4.000 ;
    END
  END out[40]
  PIN out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 421.640 4.000 422.240 ;
    END
  END out[41]
  PIN out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 880.640 1799.000 881.240 ;
    END
  END out[42]
  PIN out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.290 1.000 998.570 4.000 ;
    END
  END out[43]
  PIN out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 1796.000 1291.590 1799.000 ;
    END
  END out[44]
  PIN out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1706.690 1796.000 1706.970 1799.000 ;
    END
  END out[45]
  PIN out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 1796.000 200.010 1799.000 ;
    END
  END out[46]
  PIN out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 1.000 270.850 4.000 ;
    END
  END out[47]
  PIN out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1033.640 1799.000 1034.240 ;
    END
  END out[48]
  PIN out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1761.430 1796.000 1761.710 1799.000 ;
    END
  END out[49]
  PIN out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1169.640 4.000 1170.240 ;
    END
  END out[4]
  PIN out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1360.040 1799.000 1360.640 ;
    END
  END out[50]
  PIN out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 533.840 1799.000 534.440 ;
    END
  END out[51]
  PIN out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 1.000 1198.210 4.000 ;
    END
  END out[52]
  PIN out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.690 1796.000 1545.970 1799.000 ;
    END
  END out[53]
  PIN out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 1796.000 528.450 1799.000 ;
    END
  END out[54]
  PIN out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 1.000 544.550 4.000 ;
    END
  END out[55]
  PIN out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1050.640 1799.000 1051.240 ;
    END
  END out[56]
  PIN out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.890 1.000 1417.170 4.000 ;
    END
  END out[57]
  PIN out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 476.040 1799.000 476.640 ;
    END
  END out[58]
  PIN out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1033.640 4.000 1034.240 ;
    END
  END out[59]
  PIN out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1796.850 1.000 1797.130 4.000 ;
    END
  END out[5]
  PIN out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 1.000 290.170 4.000 ;
    END
  END out[60]
  PIN out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 1.000 853.670 4.000 ;
    END
  END out[61]
  PIN out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 727.640 1799.000 728.240 ;
    END
  END out[62]
  PIN out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.630 1796.000 1471.910 1799.000 ;
    END
  END out[63]
  PIN out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1587.840 1799.000 1588.440 ;
    END
  END out[64]
  PIN out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 34.040 1799.000 34.640 ;
    END
  END out[65]
  PIN out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 1.000 145.270 4.000 ;
    END
  END out[66]
  PIN out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 996.240 1799.000 996.840 ;
    END
  END out[67]
  PIN out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 1.000 35.790 4.000 ;
    END
  END out[68]
  PIN out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1628.640 1799.000 1629.240 ;
    END
  END out[69]
  PIN out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.570 1796.000 1397.850 1799.000 ;
    END
  END out[6]
  PIN out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 149.640 1799.000 150.240 ;
    END
  END out[70]
  PIN out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 1796.000 1327.010 1799.000 ;
    END
  END out[71]
  PIN out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 554.240 4.000 554.840 ;
    END
  END out[72]
  PIN out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 612.040 4.000 612.640 ;
    END
  END out[73]
  PIN out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.610 1.000 1178.890 4.000 ;
    END
  END out[74]
  PIN out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 1.000 0.370 4.000 ;
    END
  END out[75]
  PIN out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.250 1.000 1378.530 4.000 ;
    END
  END out[76]
  PIN out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 918.040 4.000 918.640 ;
    END
  END out[77]
  PIN out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1628.640 4.000 1629.240 ;
    END
  END out[78]
  PIN out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 1796.000 544.550 1799.000 ;
    END
  END out[79]
  PIN out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 632.440 4.000 633.040 ;
    END
  END out[7]
  PIN out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 1.000 361.010 4.000 ;
    END
  END out[80]
  PIN out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 1.000 125.950 4.000 ;
    END
  END out[81]
  PIN out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.190 1796.000 982.470 1799.000 ;
    END
  END out[82]
  PIN out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 1796.000 579.970 1799.000 ;
    END
  END out[83]
  PIN out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 1.000 943.830 4.000 ;
    END
  END out[84]
  PIN out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.990 1796.000 1272.270 1799.000 ;
    END
  END out[85]
  PIN out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 459.040 1799.000 459.640 ;
    END
  END out[86]
  PIN out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1227.440 4.000 1228.040 ;
    END
  END out[87]
  PIN out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1377.040 1799.000 1377.640 ;
    END
  END out[88]
  PIN out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 1.000 380.330 4.000 ;
    END
  END out[89]
  PIN out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 1.000 670.130 4.000 ;
    END
  END out[8]
  PIN out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 170.040 4.000 170.640 ;
    END
  END out[90]
  PIN out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1319.240 1799.000 1319.840 ;
    END
  END out[91]
  PIN out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.030 1.000 1053.310 4.000 ;
    END
  END out[92]
  PIN out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 1796.000 1198.210 1799.000 ;
    END
  END out[93]
  PIN out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.830 1796.000 1182.110 1799.000 ;
    END
  END out[94]
  PIN out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1706.840 4.000 1707.440 ;
    END
  END out[95]
  PIN out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 1796.000 235.430 1799.000 ;
    END
  END out[96]
  PIN out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.770 1.000 1269.050 4.000 ;
    END
  END out[97]
  PIN out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 401.240 4.000 401.840 ;
    END
  END out[98]
  PIN out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1533.440 4.000 1534.040 ;
    END
  END out[99]
  PIN out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 860.240 1799.000 860.840 ;
    END
  END out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 1787.280 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 1787.280 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1794.460 1787.125 ;
      LAYER met1 ;
        RECT 0.070 9.560 1797.150 1787.280 ;
      LAYER met2 ;
        RECT 0.650 1795.720 19.130 1796.290 ;
        RECT 19.970 1795.720 35.230 1796.290 ;
        RECT 36.070 1795.720 54.550 1796.290 ;
        RECT 55.390 1795.720 70.650 1796.290 ;
        RECT 71.490 1795.720 89.970 1796.290 ;
        RECT 90.810 1795.720 109.290 1796.290 ;
        RECT 110.130 1795.720 125.390 1796.290 ;
        RECT 126.230 1795.720 144.710 1796.290 ;
        RECT 145.550 1795.720 164.030 1796.290 ;
        RECT 164.870 1795.720 180.130 1796.290 ;
        RECT 180.970 1795.720 199.450 1796.290 ;
        RECT 200.290 1795.720 218.770 1796.290 ;
        RECT 219.610 1795.720 234.870 1796.290 ;
        RECT 235.710 1795.720 254.190 1796.290 ;
        RECT 255.030 1795.720 273.510 1796.290 ;
        RECT 274.350 1795.720 289.610 1796.290 ;
        RECT 290.450 1795.720 308.930 1796.290 ;
        RECT 309.770 1795.720 325.030 1796.290 ;
        RECT 325.870 1795.720 344.350 1796.290 ;
        RECT 345.190 1795.720 363.670 1796.290 ;
        RECT 364.510 1795.720 379.770 1796.290 ;
        RECT 380.610 1795.720 399.090 1796.290 ;
        RECT 399.930 1795.720 418.410 1796.290 ;
        RECT 419.250 1795.720 434.510 1796.290 ;
        RECT 435.350 1795.720 453.830 1796.290 ;
        RECT 454.670 1795.720 473.150 1796.290 ;
        RECT 473.990 1795.720 489.250 1796.290 ;
        RECT 490.090 1795.720 508.570 1796.290 ;
        RECT 509.410 1795.720 527.890 1796.290 ;
        RECT 528.730 1795.720 543.990 1796.290 ;
        RECT 544.830 1795.720 563.310 1796.290 ;
        RECT 564.150 1795.720 579.410 1796.290 ;
        RECT 580.250 1795.720 598.730 1796.290 ;
        RECT 599.570 1795.720 618.050 1796.290 ;
        RECT 618.890 1795.720 634.150 1796.290 ;
        RECT 634.990 1795.720 653.470 1796.290 ;
        RECT 654.310 1795.720 672.790 1796.290 ;
        RECT 673.630 1795.720 688.890 1796.290 ;
        RECT 689.730 1795.720 708.210 1796.290 ;
        RECT 709.050 1795.720 727.530 1796.290 ;
        RECT 728.370 1795.720 743.630 1796.290 ;
        RECT 744.470 1795.720 762.950 1796.290 ;
        RECT 763.790 1795.720 782.270 1796.290 ;
        RECT 783.110 1795.720 798.370 1796.290 ;
        RECT 799.210 1795.720 817.690 1796.290 ;
        RECT 818.530 1795.720 833.790 1796.290 ;
        RECT 834.630 1795.720 853.110 1796.290 ;
        RECT 853.950 1795.720 872.430 1796.290 ;
        RECT 873.270 1795.720 888.530 1796.290 ;
        RECT 889.370 1795.720 907.850 1796.290 ;
        RECT 908.690 1795.720 927.170 1796.290 ;
        RECT 928.010 1795.720 943.270 1796.290 ;
        RECT 944.110 1795.720 962.590 1796.290 ;
        RECT 963.430 1795.720 981.910 1796.290 ;
        RECT 982.750 1795.720 998.010 1796.290 ;
        RECT 998.850 1795.720 1017.330 1796.290 ;
        RECT 1018.170 1795.720 1036.650 1796.290 ;
        RECT 1037.490 1795.720 1052.750 1796.290 ;
        RECT 1053.590 1795.720 1072.070 1796.290 ;
        RECT 1072.910 1795.720 1088.170 1796.290 ;
        RECT 1089.010 1795.720 1107.490 1796.290 ;
        RECT 1108.330 1795.720 1126.810 1796.290 ;
        RECT 1127.650 1795.720 1142.910 1796.290 ;
        RECT 1143.750 1795.720 1162.230 1796.290 ;
        RECT 1163.070 1795.720 1181.550 1796.290 ;
        RECT 1182.390 1795.720 1197.650 1796.290 ;
        RECT 1198.490 1795.720 1216.970 1796.290 ;
        RECT 1217.810 1795.720 1236.290 1796.290 ;
        RECT 1237.130 1795.720 1252.390 1796.290 ;
        RECT 1253.230 1795.720 1271.710 1796.290 ;
        RECT 1272.550 1795.720 1291.030 1796.290 ;
        RECT 1291.870 1795.720 1307.130 1796.290 ;
        RECT 1307.970 1795.720 1326.450 1796.290 ;
        RECT 1327.290 1795.720 1342.550 1796.290 ;
        RECT 1343.390 1795.720 1361.870 1796.290 ;
        RECT 1362.710 1795.720 1381.190 1796.290 ;
        RECT 1382.030 1795.720 1397.290 1796.290 ;
        RECT 1398.130 1795.720 1416.610 1796.290 ;
        RECT 1417.450 1795.720 1435.930 1796.290 ;
        RECT 1436.770 1795.720 1452.030 1796.290 ;
        RECT 1452.870 1795.720 1471.350 1796.290 ;
        RECT 1472.190 1795.720 1490.670 1796.290 ;
        RECT 1491.510 1795.720 1506.770 1796.290 ;
        RECT 1507.610 1795.720 1526.090 1796.290 ;
        RECT 1526.930 1795.720 1545.410 1796.290 ;
        RECT 1546.250 1795.720 1561.510 1796.290 ;
        RECT 1562.350 1795.720 1580.830 1796.290 ;
        RECT 1581.670 1795.720 1596.930 1796.290 ;
        RECT 1597.770 1795.720 1616.250 1796.290 ;
        RECT 1617.090 1795.720 1635.570 1796.290 ;
        RECT 1636.410 1795.720 1651.670 1796.290 ;
        RECT 1652.510 1795.720 1670.990 1796.290 ;
        RECT 1671.830 1795.720 1690.310 1796.290 ;
        RECT 1691.150 1795.720 1706.410 1796.290 ;
        RECT 1707.250 1795.720 1725.730 1796.290 ;
        RECT 1726.570 1795.720 1745.050 1796.290 ;
        RECT 1745.890 1795.720 1761.150 1796.290 ;
        RECT 1761.990 1795.720 1780.470 1796.290 ;
        RECT 1781.310 1795.720 1796.570 1796.290 ;
        RECT 0.100 4.280 1797.120 1795.720 ;
        RECT 0.650 3.670 15.910 4.280 ;
        RECT 16.750 3.670 35.230 4.280 ;
        RECT 36.070 3.670 51.330 4.280 ;
        RECT 52.170 3.670 70.650 4.280 ;
        RECT 71.490 3.670 89.970 4.280 ;
        RECT 90.810 3.670 106.070 4.280 ;
        RECT 106.910 3.670 125.390 4.280 ;
        RECT 126.230 3.670 144.710 4.280 ;
        RECT 145.550 3.670 160.810 4.280 ;
        RECT 161.650 3.670 180.130 4.280 ;
        RECT 180.970 3.670 199.450 4.280 ;
        RECT 200.290 3.670 215.550 4.280 ;
        RECT 216.390 3.670 234.870 4.280 ;
        RECT 235.710 3.670 250.970 4.280 ;
        RECT 251.810 3.670 270.290 4.280 ;
        RECT 271.130 3.670 289.610 4.280 ;
        RECT 290.450 3.670 305.710 4.280 ;
        RECT 306.550 3.670 325.030 4.280 ;
        RECT 325.870 3.670 344.350 4.280 ;
        RECT 345.190 3.670 360.450 4.280 ;
        RECT 361.290 3.670 379.770 4.280 ;
        RECT 380.610 3.670 399.090 4.280 ;
        RECT 399.930 3.670 415.190 4.280 ;
        RECT 416.030 3.670 434.510 4.280 ;
        RECT 435.350 3.670 453.830 4.280 ;
        RECT 454.670 3.670 469.930 4.280 ;
        RECT 470.770 3.670 489.250 4.280 ;
        RECT 490.090 3.670 505.350 4.280 ;
        RECT 506.190 3.670 524.670 4.280 ;
        RECT 525.510 3.670 543.990 4.280 ;
        RECT 544.830 3.670 560.090 4.280 ;
        RECT 560.930 3.670 579.410 4.280 ;
        RECT 580.250 3.670 598.730 4.280 ;
        RECT 599.570 3.670 614.830 4.280 ;
        RECT 615.670 3.670 634.150 4.280 ;
        RECT 634.990 3.670 653.470 4.280 ;
        RECT 654.310 3.670 669.570 4.280 ;
        RECT 670.410 3.670 688.890 4.280 ;
        RECT 689.730 3.670 708.210 4.280 ;
        RECT 709.050 3.670 724.310 4.280 ;
        RECT 725.150 3.670 743.630 4.280 ;
        RECT 744.470 3.670 759.730 4.280 ;
        RECT 760.570 3.670 779.050 4.280 ;
        RECT 779.890 3.670 798.370 4.280 ;
        RECT 799.210 3.670 814.470 4.280 ;
        RECT 815.310 3.670 833.790 4.280 ;
        RECT 834.630 3.670 853.110 4.280 ;
        RECT 853.950 3.670 869.210 4.280 ;
        RECT 870.050 3.670 888.530 4.280 ;
        RECT 889.370 3.670 907.850 4.280 ;
        RECT 908.690 3.670 923.950 4.280 ;
        RECT 924.790 3.670 943.270 4.280 ;
        RECT 944.110 3.670 962.590 4.280 ;
        RECT 963.430 3.670 978.690 4.280 ;
        RECT 979.530 3.670 998.010 4.280 ;
        RECT 998.850 3.670 1014.110 4.280 ;
        RECT 1014.950 3.670 1033.430 4.280 ;
        RECT 1034.270 3.670 1052.750 4.280 ;
        RECT 1053.590 3.670 1068.850 4.280 ;
        RECT 1069.690 3.670 1088.170 4.280 ;
        RECT 1089.010 3.670 1107.490 4.280 ;
        RECT 1108.330 3.670 1123.590 4.280 ;
        RECT 1124.430 3.670 1142.910 4.280 ;
        RECT 1143.750 3.670 1162.230 4.280 ;
        RECT 1163.070 3.670 1178.330 4.280 ;
        RECT 1179.170 3.670 1197.650 4.280 ;
        RECT 1198.490 3.670 1216.970 4.280 ;
        RECT 1217.810 3.670 1233.070 4.280 ;
        RECT 1233.910 3.670 1252.390 4.280 ;
        RECT 1253.230 3.670 1268.490 4.280 ;
        RECT 1269.330 3.670 1287.810 4.280 ;
        RECT 1288.650 3.670 1307.130 4.280 ;
        RECT 1307.970 3.670 1323.230 4.280 ;
        RECT 1324.070 3.670 1342.550 4.280 ;
        RECT 1343.390 3.670 1361.870 4.280 ;
        RECT 1362.710 3.670 1377.970 4.280 ;
        RECT 1378.810 3.670 1397.290 4.280 ;
        RECT 1398.130 3.670 1416.610 4.280 ;
        RECT 1417.450 3.670 1432.710 4.280 ;
        RECT 1433.550 3.670 1452.030 4.280 ;
        RECT 1452.870 3.670 1471.350 4.280 ;
        RECT 1472.190 3.670 1487.450 4.280 ;
        RECT 1488.290 3.670 1506.770 4.280 ;
        RECT 1507.610 3.670 1522.870 4.280 ;
        RECT 1523.710 3.670 1542.190 4.280 ;
        RECT 1543.030 3.670 1561.510 4.280 ;
        RECT 1562.350 3.670 1577.610 4.280 ;
        RECT 1578.450 3.670 1596.930 4.280 ;
        RECT 1597.770 3.670 1616.250 4.280 ;
        RECT 1617.090 3.670 1632.350 4.280 ;
        RECT 1633.190 3.670 1651.670 4.280 ;
        RECT 1652.510 3.670 1670.990 4.280 ;
        RECT 1671.830 3.670 1687.090 4.280 ;
        RECT 1687.930 3.670 1706.410 4.280 ;
        RECT 1707.250 3.670 1725.730 4.280 ;
        RECT 1726.570 3.670 1741.830 4.280 ;
        RECT 1742.670 3.670 1761.150 4.280 ;
        RECT 1761.990 3.670 1777.250 4.280 ;
        RECT 1778.090 3.670 1796.570 4.280 ;
      LAYER met3 ;
        RECT 4.000 1782.640 1796.000 1787.205 ;
        RECT 4.400 1781.240 1795.600 1782.640 ;
        RECT 4.000 1765.640 1796.000 1781.240 ;
        RECT 4.400 1764.240 1796.000 1765.640 ;
        RECT 4.000 1762.240 1796.000 1764.240 ;
        RECT 4.000 1760.840 1795.600 1762.240 ;
        RECT 4.000 1745.240 1796.000 1760.840 ;
        RECT 4.400 1743.840 1795.600 1745.240 ;
        RECT 4.000 1724.840 1796.000 1743.840 ;
        RECT 4.400 1723.440 1795.600 1724.840 ;
        RECT 4.000 1707.840 1796.000 1723.440 ;
        RECT 4.400 1706.440 1796.000 1707.840 ;
        RECT 4.000 1704.440 1796.000 1706.440 ;
        RECT 4.000 1703.040 1795.600 1704.440 ;
        RECT 4.000 1687.440 1796.000 1703.040 ;
        RECT 4.400 1686.040 1795.600 1687.440 ;
        RECT 4.000 1667.040 1796.000 1686.040 ;
        RECT 4.400 1665.640 1795.600 1667.040 ;
        RECT 4.000 1650.040 1796.000 1665.640 ;
        RECT 4.400 1648.640 1796.000 1650.040 ;
        RECT 4.000 1646.640 1796.000 1648.640 ;
        RECT 4.000 1645.240 1795.600 1646.640 ;
        RECT 4.000 1629.640 1796.000 1645.240 ;
        RECT 4.400 1628.240 1795.600 1629.640 ;
        RECT 4.000 1609.240 1796.000 1628.240 ;
        RECT 4.400 1607.840 1795.600 1609.240 ;
        RECT 4.000 1592.240 1796.000 1607.840 ;
        RECT 4.400 1590.840 1796.000 1592.240 ;
        RECT 4.000 1588.840 1796.000 1590.840 ;
        RECT 4.000 1587.440 1795.600 1588.840 ;
        RECT 4.000 1571.840 1796.000 1587.440 ;
        RECT 4.400 1570.440 1795.600 1571.840 ;
        RECT 4.000 1554.840 1796.000 1570.440 ;
        RECT 4.400 1553.440 1796.000 1554.840 ;
        RECT 4.000 1551.440 1796.000 1553.440 ;
        RECT 4.000 1550.040 1795.600 1551.440 ;
        RECT 4.000 1534.440 1796.000 1550.040 ;
        RECT 4.400 1533.040 1795.600 1534.440 ;
        RECT 4.000 1514.040 1796.000 1533.040 ;
        RECT 4.400 1512.640 1795.600 1514.040 ;
        RECT 4.000 1497.040 1796.000 1512.640 ;
        RECT 4.400 1495.640 1796.000 1497.040 ;
        RECT 4.000 1493.640 1796.000 1495.640 ;
        RECT 4.000 1492.240 1795.600 1493.640 ;
        RECT 4.000 1476.640 1796.000 1492.240 ;
        RECT 4.400 1475.240 1795.600 1476.640 ;
        RECT 4.000 1456.240 1796.000 1475.240 ;
        RECT 4.400 1454.840 1795.600 1456.240 ;
        RECT 4.000 1439.240 1796.000 1454.840 ;
        RECT 4.400 1437.840 1796.000 1439.240 ;
        RECT 4.000 1435.840 1796.000 1437.840 ;
        RECT 4.000 1434.440 1795.600 1435.840 ;
        RECT 4.000 1418.840 1796.000 1434.440 ;
        RECT 4.400 1417.440 1795.600 1418.840 ;
        RECT 4.000 1398.440 1796.000 1417.440 ;
        RECT 4.400 1397.040 1795.600 1398.440 ;
        RECT 4.000 1381.440 1796.000 1397.040 ;
        RECT 4.400 1380.040 1796.000 1381.440 ;
        RECT 4.000 1378.040 1796.000 1380.040 ;
        RECT 4.000 1376.640 1795.600 1378.040 ;
        RECT 4.000 1361.040 1796.000 1376.640 ;
        RECT 4.400 1359.640 1795.600 1361.040 ;
        RECT 4.000 1340.640 1796.000 1359.640 ;
        RECT 4.400 1339.240 1795.600 1340.640 ;
        RECT 4.000 1323.640 1796.000 1339.240 ;
        RECT 4.400 1322.240 1796.000 1323.640 ;
        RECT 4.000 1320.240 1796.000 1322.240 ;
        RECT 4.000 1318.840 1795.600 1320.240 ;
        RECT 4.000 1303.240 1796.000 1318.840 ;
        RECT 4.400 1301.840 1795.600 1303.240 ;
        RECT 4.000 1286.240 1796.000 1301.840 ;
        RECT 4.400 1284.840 1796.000 1286.240 ;
        RECT 4.000 1282.840 1796.000 1284.840 ;
        RECT 4.000 1281.440 1795.600 1282.840 ;
        RECT 4.000 1265.840 1796.000 1281.440 ;
        RECT 4.400 1264.440 1795.600 1265.840 ;
        RECT 4.000 1245.440 1796.000 1264.440 ;
        RECT 4.400 1244.040 1795.600 1245.440 ;
        RECT 4.000 1228.440 1796.000 1244.040 ;
        RECT 4.400 1227.040 1796.000 1228.440 ;
        RECT 4.000 1225.040 1796.000 1227.040 ;
        RECT 4.000 1223.640 1795.600 1225.040 ;
        RECT 4.000 1208.040 1796.000 1223.640 ;
        RECT 4.400 1206.640 1795.600 1208.040 ;
        RECT 4.000 1187.640 1796.000 1206.640 ;
        RECT 4.400 1186.240 1795.600 1187.640 ;
        RECT 4.000 1170.640 1796.000 1186.240 ;
        RECT 4.400 1169.240 1796.000 1170.640 ;
        RECT 4.000 1167.240 1796.000 1169.240 ;
        RECT 4.000 1165.840 1795.600 1167.240 ;
        RECT 4.000 1150.240 1796.000 1165.840 ;
        RECT 4.400 1148.840 1795.600 1150.240 ;
        RECT 4.000 1129.840 1796.000 1148.840 ;
        RECT 4.400 1128.440 1795.600 1129.840 ;
        RECT 4.000 1112.840 1796.000 1128.440 ;
        RECT 4.400 1111.440 1796.000 1112.840 ;
        RECT 4.000 1109.440 1796.000 1111.440 ;
        RECT 4.000 1108.040 1795.600 1109.440 ;
        RECT 4.000 1092.440 1796.000 1108.040 ;
        RECT 4.400 1091.040 1795.600 1092.440 ;
        RECT 4.000 1072.040 1796.000 1091.040 ;
        RECT 4.400 1070.640 1795.600 1072.040 ;
        RECT 4.000 1055.040 1796.000 1070.640 ;
        RECT 4.400 1053.640 1796.000 1055.040 ;
        RECT 4.000 1051.640 1796.000 1053.640 ;
        RECT 4.000 1050.240 1795.600 1051.640 ;
        RECT 4.000 1034.640 1796.000 1050.240 ;
        RECT 4.400 1033.240 1795.600 1034.640 ;
        RECT 4.000 1017.640 1796.000 1033.240 ;
        RECT 4.400 1016.240 1796.000 1017.640 ;
        RECT 4.000 1014.240 1796.000 1016.240 ;
        RECT 4.000 1012.840 1795.600 1014.240 ;
        RECT 4.000 997.240 1796.000 1012.840 ;
        RECT 4.400 995.840 1795.600 997.240 ;
        RECT 4.000 976.840 1796.000 995.840 ;
        RECT 4.400 975.440 1795.600 976.840 ;
        RECT 4.000 959.840 1796.000 975.440 ;
        RECT 4.400 958.440 1796.000 959.840 ;
        RECT 4.000 956.440 1796.000 958.440 ;
        RECT 4.000 955.040 1795.600 956.440 ;
        RECT 4.000 939.440 1796.000 955.040 ;
        RECT 4.400 938.040 1795.600 939.440 ;
        RECT 4.000 919.040 1796.000 938.040 ;
        RECT 4.400 917.640 1795.600 919.040 ;
        RECT 4.000 902.040 1796.000 917.640 ;
        RECT 4.400 900.640 1796.000 902.040 ;
        RECT 4.000 898.640 1796.000 900.640 ;
        RECT 4.000 897.240 1795.600 898.640 ;
        RECT 4.000 881.640 1796.000 897.240 ;
        RECT 4.400 880.240 1795.600 881.640 ;
        RECT 4.000 861.240 1796.000 880.240 ;
        RECT 4.400 859.840 1795.600 861.240 ;
        RECT 4.000 844.240 1796.000 859.840 ;
        RECT 4.400 842.840 1796.000 844.240 ;
        RECT 4.000 840.840 1796.000 842.840 ;
        RECT 4.000 839.440 1795.600 840.840 ;
        RECT 4.000 823.840 1796.000 839.440 ;
        RECT 4.400 822.440 1795.600 823.840 ;
        RECT 4.000 803.440 1796.000 822.440 ;
        RECT 4.400 802.040 1795.600 803.440 ;
        RECT 4.000 786.440 1796.000 802.040 ;
        RECT 4.400 785.040 1796.000 786.440 ;
        RECT 4.000 783.040 1796.000 785.040 ;
        RECT 4.000 781.640 1795.600 783.040 ;
        RECT 4.000 766.040 1796.000 781.640 ;
        RECT 4.400 764.640 1795.600 766.040 ;
        RECT 4.000 749.040 1796.000 764.640 ;
        RECT 4.400 747.640 1796.000 749.040 ;
        RECT 4.000 745.640 1796.000 747.640 ;
        RECT 4.000 744.240 1795.600 745.640 ;
        RECT 4.000 728.640 1796.000 744.240 ;
        RECT 4.400 727.240 1795.600 728.640 ;
        RECT 4.000 708.240 1796.000 727.240 ;
        RECT 4.400 706.840 1795.600 708.240 ;
        RECT 4.000 691.240 1796.000 706.840 ;
        RECT 4.400 689.840 1796.000 691.240 ;
        RECT 4.000 687.840 1796.000 689.840 ;
        RECT 4.000 686.440 1795.600 687.840 ;
        RECT 4.000 670.840 1796.000 686.440 ;
        RECT 4.400 669.440 1795.600 670.840 ;
        RECT 4.000 650.440 1796.000 669.440 ;
        RECT 4.400 649.040 1795.600 650.440 ;
        RECT 4.000 633.440 1796.000 649.040 ;
        RECT 4.400 632.040 1796.000 633.440 ;
        RECT 4.000 630.040 1796.000 632.040 ;
        RECT 4.000 628.640 1795.600 630.040 ;
        RECT 4.000 613.040 1796.000 628.640 ;
        RECT 4.400 611.640 1795.600 613.040 ;
        RECT 4.000 592.640 1796.000 611.640 ;
        RECT 4.400 591.240 1795.600 592.640 ;
        RECT 4.000 575.640 1796.000 591.240 ;
        RECT 4.400 574.240 1796.000 575.640 ;
        RECT 4.000 572.240 1796.000 574.240 ;
        RECT 4.000 570.840 1795.600 572.240 ;
        RECT 4.000 555.240 1796.000 570.840 ;
        RECT 4.400 553.840 1795.600 555.240 ;
        RECT 4.000 534.840 1796.000 553.840 ;
        RECT 4.400 533.440 1795.600 534.840 ;
        RECT 4.000 517.840 1796.000 533.440 ;
        RECT 4.400 516.440 1796.000 517.840 ;
        RECT 4.000 514.440 1796.000 516.440 ;
        RECT 4.000 513.040 1795.600 514.440 ;
        RECT 4.000 497.440 1796.000 513.040 ;
        RECT 4.400 496.040 1795.600 497.440 ;
        RECT 4.000 480.440 1796.000 496.040 ;
        RECT 4.400 479.040 1796.000 480.440 ;
        RECT 4.000 477.040 1796.000 479.040 ;
        RECT 4.000 475.640 1795.600 477.040 ;
        RECT 4.000 460.040 1796.000 475.640 ;
        RECT 4.400 458.640 1795.600 460.040 ;
        RECT 4.000 439.640 1796.000 458.640 ;
        RECT 4.400 438.240 1795.600 439.640 ;
        RECT 4.000 422.640 1796.000 438.240 ;
        RECT 4.400 421.240 1796.000 422.640 ;
        RECT 4.000 419.240 1796.000 421.240 ;
        RECT 4.000 417.840 1795.600 419.240 ;
        RECT 4.000 402.240 1796.000 417.840 ;
        RECT 4.400 400.840 1795.600 402.240 ;
        RECT 4.000 381.840 1796.000 400.840 ;
        RECT 4.400 380.440 1795.600 381.840 ;
        RECT 4.000 364.840 1796.000 380.440 ;
        RECT 4.400 363.440 1796.000 364.840 ;
        RECT 4.000 361.440 1796.000 363.440 ;
        RECT 4.000 360.040 1795.600 361.440 ;
        RECT 4.000 344.440 1796.000 360.040 ;
        RECT 4.400 343.040 1795.600 344.440 ;
        RECT 4.000 324.040 1796.000 343.040 ;
        RECT 4.400 322.640 1795.600 324.040 ;
        RECT 4.000 307.040 1796.000 322.640 ;
        RECT 4.400 305.640 1796.000 307.040 ;
        RECT 4.000 303.640 1796.000 305.640 ;
        RECT 4.000 302.240 1795.600 303.640 ;
        RECT 4.000 286.640 1796.000 302.240 ;
        RECT 4.400 285.240 1795.600 286.640 ;
        RECT 4.000 266.240 1796.000 285.240 ;
        RECT 4.400 264.840 1795.600 266.240 ;
        RECT 4.000 249.240 1796.000 264.840 ;
        RECT 4.400 247.840 1796.000 249.240 ;
        RECT 4.000 245.840 1796.000 247.840 ;
        RECT 4.000 244.440 1795.600 245.840 ;
        RECT 4.000 228.840 1796.000 244.440 ;
        RECT 4.400 227.440 1795.600 228.840 ;
        RECT 4.000 211.840 1796.000 227.440 ;
        RECT 4.400 210.440 1796.000 211.840 ;
        RECT 4.000 208.440 1796.000 210.440 ;
        RECT 4.000 207.040 1795.600 208.440 ;
        RECT 4.000 191.440 1796.000 207.040 ;
        RECT 4.400 190.040 1795.600 191.440 ;
        RECT 4.000 171.040 1796.000 190.040 ;
        RECT 4.400 169.640 1795.600 171.040 ;
        RECT 4.000 154.040 1796.000 169.640 ;
        RECT 4.400 152.640 1796.000 154.040 ;
        RECT 4.000 150.640 1796.000 152.640 ;
        RECT 4.000 149.240 1795.600 150.640 ;
        RECT 4.000 133.640 1796.000 149.240 ;
        RECT 4.400 132.240 1795.600 133.640 ;
        RECT 4.000 113.240 1796.000 132.240 ;
        RECT 4.400 111.840 1795.600 113.240 ;
        RECT 4.000 96.240 1796.000 111.840 ;
        RECT 4.400 94.840 1796.000 96.240 ;
        RECT 4.000 92.840 1796.000 94.840 ;
        RECT 4.000 91.440 1795.600 92.840 ;
        RECT 4.000 75.840 1796.000 91.440 ;
        RECT 4.400 74.440 1795.600 75.840 ;
        RECT 4.000 55.440 1796.000 74.440 ;
        RECT 4.400 54.040 1795.600 55.440 ;
        RECT 4.000 38.440 1796.000 54.040 ;
        RECT 4.400 37.040 1796.000 38.440 ;
        RECT 4.000 35.040 1796.000 37.040 ;
        RECT 4.000 33.640 1795.600 35.040 ;
        RECT 4.000 18.040 1796.000 33.640 ;
        RECT 4.400 16.640 1795.600 18.040 ;
        RECT 4.000 7.655 1796.000 16.640 ;
      LAYER met4 ;
        RECT 31.575 10.240 97.440 1786.185 ;
        RECT 99.840 10.240 174.240 1786.185 ;
        RECT 176.640 10.240 251.040 1786.185 ;
        RECT 253.440 10.240 327.840 1786.185 ;
        RECT 330.240 10.240 404.640 1786.185 ;
        RECT 407.040 10.240 481.440 1786.185 ;
        RECT 483.840 10.240 558.240 1786.185 ;
        RECT 560.640 10.240 635.040 1786.185 ;
        RECT 637.440 10.240 711.840 1786.185 ;
        RECT 714.240 10.240 788.640 1786.185 ;
        RECT 791.040 10.240 865.440 1786.185 ;
        RECT 867.840 10.240 942.240 1786.185 ;
        RECT 944.640 10.240 1019.040 1786.185 ;
        RECT 1021.440 10.240 1095.840 1786.185 ;
        RECT 1098.240 10.240 1172.640 1786.185 ;
        RECT 1175.040 10.240 1249.440 1786.185 ;
        RECT 1251.840 10.240 1326.240 1786.185 ;
        RECT 1328.640 10.240 1403.040 1786.185 ;
        RECT 1405.440 10.240 1479.840 1786.185 ;
        RECT 1482.240 10.240 1556.640 1786.185 ;
        RECT 1559.040 10.240 1633.440 1786.185 ;
        RECT 1635.840 10.240 1710.240 1786.185 ;
        RECT 1712.640 10.240 1768.865 1786.185 ;
        RECT 31.575 7.655 1768.865 10.240 ;
  END
END decrypt_aes128
END LIBRARY

